module medium_1 ( clock, 
    n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, n3070gat, n3071gat,
    n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, n3077gat, n3078gat,
    n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, n3084gat, n3085gat,
    n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat, n3092gat,
    n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, n3099gat, n3100gat,
    n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat,
    n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat,
    n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat,
    n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat,
    n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat,
    n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat,
    n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat  );
  input  clock, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, n3070gat,
    n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, n3077gat,
    n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, n3084gat,
    n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat,
    n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, n3099gat,
    n3100gat;
  output n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat,
    n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat,
    n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat,
    n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat,
    n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat,
    n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat,
    n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat;
  reg n673gat, n398gat, n402gat, n919gat, n846gat, n394gat, n703gat,
    n722gat, n726gat, n2510gat, n271gat, n160gat, n337gat, n842gat,
    n341gat, n2522gat, n2472gat, n2319gat, n1821gat, n1825gat, n2029gat,
    n1829gat, n283gat, n165gat, n279gat, n1026gat, n275gat, n2476gat,
    n1068gat, n957gat, n861gat, n1294gat, n1241gat, n1298gat, n865gat,
    n1080gat, n1148gat, n2468gat, n618gat, n491gat, n622gat, n626gat,
    n834gat, n707gat, n838gat, n830gat, n614gat, n2526gat, n680gat,
    n816gat, n580gat, n824gat, n820gat, n883gat, n584gat, n684gat, n699gat,
    n2464gat, n2399gat, n2343gat, n2203gat, n2562gat, n2207gat, n2626gat,
    n2490gat, n2622gat, n2630gat, n2543gat, n2102gat, n1880gat, n1763gat,
    n2155gat, n1035gat, n1121gat, n1072gat, n1282gat, n1226gat, n931gat,
    n1135gat, n1045gat, n1197gat, n2518gat, n667gat, n659gat, n553gat,
    n777gat, n561gat, n366gat, n322gat, n318gat, n314gat, n2599gat,
    n2588gat, n2640gat, n2658gat, n2495gat, n2390gat, n2270gat, n2339gat,
    n2502gat, n2634gat, n2506gat, n1834gat, n1767gat, n2084gat, n2143gat,
    n2061gat, n2139gat, n1899gat, n1850gat, n2403gat, n2394gat, n2440gat,
    n2407gat, n2347gat, n1389gat, n2021gat, n1394gat, n1496gat, n2091gat,
    n1332gat, n1740gat, n2179gat, n2190gat, n2135gat, n2262gat, n2182gat,
    n1433gat, n1316gat, n1363gat, n1312gat, n1775gat, n1871gat, n2592gat,
    n1508gat, n1678gat, n2309gat, n2450gat, n2446gat, n2095gat, n2176gat,
    n2169gat, n2454gat, n2040gat, n2044gat, n2037gat, n2025gat, n2099gat,
    n2266gat, n2033gat, n2110gat, n2125gat, n2121gat, n2117gat, n1975gat,
    n2644gat, n156gat, n152gat, n331gat, n388gat, n463gat, n327gat,
    n384gat, n256gat, n470gat, n148gat, n2458gat, n2514gat, n1771gat,
    n1336gat, n1748gat, n1675gat, n1807gat, n1340gat, n1456gat, n1525gat,
    n1462gat, n1596gat, n1588gat;
  wire n623, n624_1, n625, n626, n627, n628, n629_1, n630, n631, n632, n633,
    n634_1, n635, n636, n637, n638, n640, n641, n642, n643, n644_1, n645,
    n646, n647, n649_1, n651, n652, n653, n654_1, n655, n657, n658, n659_1,
    n660, n662, n663, n664_1, n666, n667, n668, n670, n671, n672, n673,
    n675, n676, n677, n678, n679_1, n680, n681, n682, n683, n684_1, n685,
    n686, n687, n688, n689_1, n690, n691, n692, n693, n694_1, n695, n697,
    n698, n699_1, n700, n701, n702, n703, n704_1, n705, n706, n707, n708,
    n709_1, n710, n711, n712, n713, n714_1, n715, n716, n717, n718, n719_1,
    n720, n721, n722, n723, n724_1, n725, n726, n727, n728, n729_1, n730,
    n731, n732, n733, n734_1, n735, n736, n737, n739_1, n740, n741, n742,
    n743, n744_1, n745, n746, n747, n748, n749_1, n750, n751, n752, n753,
    n754_1, n755, n756, n757, n758, n759_1, n760, n761, n762, n763, n764_1,
    n766, n767, n768, n769_1, n770, n771, n772, n773, n774_1, n775, n776,
    n777, n778, n779_1, n780, n781, n782, n783, n784_1, n785, n786, n787,
    n788, n789_1, n790, n791, n793, n794_1, n795, n796, n797, n798, n799_1,
    n800, n801, n802, n803, n804_1, n805, n806, n807, n808, n809_1, n810,
    n811, n812, n813, n814_1, n815, n816, n817, n818, n820, n821, n822,
    n823, n824_1, n825, n826, n827, n828, n829_1, n830, n831, n832, n833,
    n834_1, n835, n836, n837, n838, n839_1, n840, n841, n842, n843, n844_1,
    n845, n847, n848, n849_1, n850, n851, n852, n853, n854_1, n855, n856,
    n857, n858, n859_1, n860, n861, n862, n863, n864_1, n865, n866, n867,
    n868, n869_1, n870, n871, n872, n874_1, n875, n876, n877, n878, n879_1,
    n880, n881, n882, n883, n884_1, n885, n886, n887, n888, n889_1, n890,
    n891, n892, n893, n894_1, n895, n896, n897, n898, n899_1, n900, n902,
    n903, n904_1, n905, n906, n907, n908, n909_1, n910, n911, n912, n914_1,
    n915, n916, n917, n918, n919_1, n920, n921, n922, n923, n924_1, n925,
    n926, n927, n928, n929_1, n931, n932, n933, n934_1, n935, n936, n937,
    n938, n939_1, n940, n941, n942, n943, n944_1, n945, n946, n947, n949_1,
    n950, n951, n952, n953, n954_1, n956, n957, n958, n959_1, n960, n961,
    n963, n964_1, n965, n966, n967, n968, n970, n971, n972, n973, n974_1,
    n975, n977, n978, n979_1, n980, n981, n982, n984_1, n985, n986, n987,
    n988, n989_1, n991, n992, n993, n994_1, n995, n996, n998, n999_1,
    n1000, n1001, n1002, n1003, n1005, n1006, n1007, n1008, n1009_1, n1010,
    n1011, n1012, n1013, n1014_1, n1015, n1016, n1017, n1018, n1019_1,
    n1020, n1021, n1022, n1023, n1024_1, n1025, n1026, n1027, n1028,
    n1029_1, n1030, n1031, n1032, n1033, n1034_1, n1035, n1036, n1037,
    n1038, n1039_1, n1040, n1041, n1042, n1043, n1044_1, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
    n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1154, n1155, n1156, n1157, n1158,
    n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1169,
    n1171, n1172, n1174, n1175, n1176, n1177, n1179, n1180, n1181, n1182,
    n1183, n1184, n1188, n1189, n1191, n1192, n1194, n1195, n1197, n1198,
    n1200, n1201, n1203, n1204, n1206, n1207, n1209, n1210, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1223, n1224,
    n1225, n1226, n1227, n1228, n1230, n1231, n1232, n1233, n1234, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1245, n1246, n1247,
    n1248, n1250, n1251, n1252, n1254, n1255, n1257, n1258, n1260, n1261,
    n1262, n1263, n1264, n1265, n1266, n1267, n1269, n1270, n1271, n1272,
    n1273, n1274, n1275, n1276, n1277, n1279, n1280, n1281, n1282, n1283,
    n1285, n1286, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1305, n1306, n1307, n1308,
    n1309, n1311, n1312, n1313, n1314, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1327, n1328, n1329, n1330, n1338, n1340, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349, n1351, n1353, n1355, n1357,
    n1359, n1361, n1363, n1365, n1367, n1368, n1369, n1370, n1372, n1373,
    n1375, n1376, n1378, n1379, n1381, n1382, n1384, n1385, n1387, n1388,
    n1390, n1391, n1393, n1394, n1397, n1398, n1399, n1400, n1402, n1403,
    n1407, n1408, n1409, n1410, n1414, n1415, n1416, n1417, n1420, n1424,
    n1425, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1451, n1452, n169, n174, n179, n184, n189, n193, n197, n201,
    n205, n210, n215, n220, n225, n230, n235, n240, n245, n250, n255, n259,
    n264, n269, n273, n277, n281, n285, n289, n294, n299, n304, n309, n314,
    n319, n323, n328, n333, n338, n343, n347, n351, n355, n359, n364, n369,
    n374, n379, n384, n389, n394, n399, n404, n409, n414, n419, n424, n429,
    n434, n439, n444, n449, n454, n459, n464, n469, n474, n479, n484, n489,
    n494, n499, n504, n509, n514, n519, n524, n529, n534, n539, n544, n549,
    n554, n559, n564, n569, n574, n579, n584, n589, n594, n599, n604, n609,
    n614, n619, n624, n629, n634, n639, n644, n649, n654, n659, n664, n669,
    n674, n679, n684, n689, n694, n699, n704, n709, n714, n719, n724, n729,
    n734, n739, n744, n749, n754, n759, n764, n769, n774, n779, n784, n789,
    n794, n799, n804, n809, n814, n819, n824, n829, n834, n839, n844, n849,
    n854, n859, n864, n869, n874, n879, n884, n889, n894, n899, n904, n909,
    n914, n919, n924, n929, n934, n939, n944, n949, n954, n959, n964, n969,
    n974, n979, n984, n989, n994, n999, n1004, n1009, n1014, n1019, n1024,
    n1029, n1034, n1039, n1044;
  assign n3112gat = 1'b1;
  assign n3104gat = n623 | ~n629_1 | n634_1;
  assign n623 = n3094gat & n624_1;
  assign n624_1 = ~n625 & n627 & ~n628;
  assign n625 = n3086gat & n626;
  assign n626 = n3095gat & ~n3083gat & ~n3085gat & ~n3084gat & n1871gat;
  assign n627 = n3087gat & n626;
  assign n628 = n3088gat & n626;
  assign n629_1 = ~n630 & ~n633;
  assign n630 = n1850gat & n631;
  assign n631 = ~n2061gat & n632 & ~n2143gat;
  assign n632 = ~n2139gat & ~n1899gat;
  assign n633 = ~n1850gat & ~n631;
  assign n634_1 = n635 & ~n638;
  assign n635 = n3086gat & ~n3085gat & n636 & n637;
  assign n636 = ~n3084gat & n1871gat & ~n3083gat & n3093gat;
  assign n637 = ~n3087gat & n3088gat;
  assign n638 = ~n3091gat & ~n3092gat;
  assign n3105gat = n640 | ~n642 | n646;
  assign n640 = ~n628 & n641 & ~n627;
  assign n641 = n3094gat & n625;
  assign n642 = ~n645 & ~n643 & ~n644_1;
  assign n643 = ~n2061gat & n632 & n2143gat;
  assign n644_1 = ~n2143gat & n2061gat;
  assign n645 = ~n2143gat & ~n632;
  assign n646 = n647 & n637 & n636 & ~n638;
  assign n647 = n3085gat & ~n3086gat;
  assign n3107gat = n1871gat & ~n649_1;
  assign n649_1 = n1775gat & n1771gat;
  assign n3108gat = ~n1035gat | ~n651;
  assign n651 = ~n652 & ~n655;
  assign n652 = n2407gat & n653;
  assign n653 = ~n2347gat & n654_1 & ~n2403gat;
  assign n654_1 = ~n2394gat & ~n2440gat;
  assign n655 = ~n2407gat & ~n653;
  assign n3109gat = ~n1072gat | ~n657;
  assign n657 = ~n660 & ~n658 & ~n659_1;
  assign n658 = ~n2347gat & ~n654_1;
  assign n659_1 = n2347gat & n654_1 & ~n2403gat;
  assign n660 = n2403gat & ~n2347gat;
  assign n3110gat = ~n1121gat | ~n662;
  assign n662 = ~n663 & ~n664_1;
  assign n663 = ~n2403gat & ~n654_1;
  assign n664_1 = n2403gat & n654_1;
  assign n3111gat = ~n931gat | ~n666;
  assign n666 = ~n667 & n2394gat & ~n668;
  assign n667 = n2394gat & ~n2440gat;
  assign n668 = ~n2394gat & n2440gat;
  assign n3113gat = ~n1135gat | ~n670;
  assign n670 = ~n671 & ~n673;
  assign n671 = n2135gat & n672;
  assign n672 = ~n2190gat & ~n2262gat;
  assign n673 = ~n2135gat & ~n672;
  assign n3114gat = ~n1282gat | ~n675;
  assign n675 = ~n676 & n2190gat & ~n677;
  assign n676 = n2190gat & ~n2262gat;
  assign n677 = ~n2190gat & n2262gat;
  assign n678 = ~n695 & ~n694_1 & ~n679_1 & ~n693;
  assign n679_1 = n690 & ~n680 & ~n685;
  assign n680 = ~n684_1 & ~n683 & ~n681 & ~n682;
  assign n681 = ~n1135gat & ~n1045gat & ~n931gat;
  assign n682 = n1135gat & n1045gat & ~n931gat;
  assign n683 = ~n1045gat & n931gat & n1135gat;
  assign n684_1 = ~n1135gat & n1045gat & n931gat;
  assign n685 = ~n689_1 & ~n688 & ~n686 & ~n687;
  assign n686 = ~n1121gat & ~n1072gat & ~n1035gat;
  assign n687 = n1121gat & n1072gat & ~n1035gat;
  assign n688 = ~n1072gat & n1035gat & n1121gat;
  assign n689_1 = ~n1121gat & n1072gat & n1035gat;
  assign n690 = ~n691 & ~n692;
  assign n691 = n1282gat & ~n1226gat;
  assign n692 = ~n1282gat & n1226gat;
  assign n693 = ~n690 & n680 & ~n685;
  assign n694_1 = ~n680 & n685 & ~n690;
  assign n695 = n690 & n680 & n685;
  assign n3117gat = n697 | n722;
  assign n697 = ~n698 & n716;
  assign n698 = ~n714_1 & ~n712 & ~n699_1 & ~n710;
  assign n699_1 = ~n271gat & n700;
  assign n700 = ~n707 & ~n701 & ~n704_1;
  assign n701 = ~n702 & ~n703;
  assign n702 = n3086gat & n3093gat;
  assign n703 = n3087gat & n3095gat;
  assign n704_1 = ~n705 & ~n706;
  assign n705 = n3087gat & n3093gat;
  assign n706 = n3088gat & n3095gat;
  assign n707 = ~n708 & ~n709_1;
  assign n708 = n3085gat & n3093gat;
  assign n709_1 = n3086gat & n3095gat;
  assign n710 = ~n1068gat & n711;
  assign n711 = n707 & ~n701 & ~n704_1;
  assign n712 = ~n680gat & n713;
  assign n713 = ~n707 & n701 & ~n704_1;
  assign n714_1 = ~n659gat & n715;
  assign n715 = ~n707 & n704_1 & ~n701;
  assign n716 = n717 & ~n721;
  assign n717 = ~n720 & ~n718 & ~n719_1;
  assign n718 = n3084gat & n3095gat;
  assign n719_1 = n3085gat & n3095gat;
  assign n720 = n3083gat & n3095gat;
  assign n721 = ~n703 & ~n709_1;
  assign n722 = ~n737 & ~n736 & ~n723 & ~n735;
  assign n723 = n732 & ~n724_1 & ~n729_1;
  assign n724_1 = ~n728 & ~n727 & ~n725 & ~n726;
  assign n725 = n3085gat & n3084gat & n3083gat;
  assign n726 = ~n3084gat & n3083gat & ~n3085gat;
  assign n727 = ~n3085gat & n3084gat & ~n3083gat;
  assign n728 = n3085gat & ~n3084gat & ~n3083gat;
  assign n729_1 = ~n730 & ~n731;
  assign n730 = n3086gat & ~n3087gat;
  assign n731 = ~n3086gat & n3087gat;
  assign n732 = ~n733 & ~n734_1;
  assign n733 = ~n3088gat & n3089gat;
  assign n734_1 = n3088gat & ~n3089gat;
  assign n735 = ~n724_1 & n729_1 & ~n732;
  assign n736 = ~n732 & n724_1 & ~n729_1;
  assign n737 = n732 & n724_1 & n729_1;
  assign n3118gat = n739_1 | n745;
  assign n739_1 = n716 & ~n740;
  assign n740 = ~n744_1 & ~n743 & ~n741 & ~n742;
  assign n741 = ~n337gat & n700;
  assign n742 = ~n861gat & n711;
  assign n743 = ~n580gat & n713;
  assign n744_1 = ~n777gat & n715;
  assign n745 = ~n764_1 & ~n763 & ~n746 & ~n762;
  assign n746 = n757 & ~n747 & ~n752;
  assign n747 = ~n751 & ~n750 & ~n748 & ~n749_1;
  assign n748 = ~n341gat & ~n394gat & ~n703gat;
  assign n749_1 = ~n341gat & n394gat & n703gat;
  assign n750 = ~n394gat & n703gat & n341gat;
  assign n751 = n341gat & n394gat & ~n703gat;
  assign n752 = ~n756 & ~n755 & ~n753 & ~n754_1;
  assign n753 = ~n160gat & ~n337gat & ~n271gat;
  assign n754_1 = n160gat & n337gat & ~n271gat;
  assign n755 = ~n337gat & n271gat & n160gat;
  assign n756 = ~n160gat & n337gat & n271gat;
  assign n757 = ~n761 & ~n760 & ~n758 & ~n759_1;
  assign n758 = ~n842gat & ~n722gat & ~n726gat;
  assign n759_1 = n842gat & n722gat & ~n726gat;
  assign n760 = ~n722gat & n726gat & n842gat;
  assign n761 = ~n842gat & n722gat & n726gat;
  assign n762 = ~n757 & n747 & ~n752;
  assign n763 = ~n747 & n752 & ~n757;
  assign n764_1 = n757 & n747 & n752;
  assign n3119gat = n766 | n772;
  assign n766 = n716 & ~n767;
  assign n767 = ~n771 & ~n770 & ~n768 & ~n769_1;
  assign n768 = ~n957gat & n711;
  assign n769_1 = ~n553gat & n715;
  assign n770 = ~n160gat & n700;
  assign n771 = ~n816gat & n713;
  assign n772 = ~n791 & ~n790 & ~n773 & ~n789_1;
  assign n773 = n784_1 & ~n774_1 & ~n779_1;
  assign n774_1 = ~n778 & ~n777 & ~n775 & ~n776;
  assign n775 = ~n1080gat & ~n1148gat & ~n865gat;
  assign n776 = n1080gat & n1148gat & ~n865gat;
  assign n777 = ~n1148gat & n865gat & n1080gat;
  assign n778 = ~n1080gat & n1148gat & n865gat;
  assign n779_1 = ~n783 & ~n782 & ~n780 & ~n781;
  assign n780 = ~n957gat & ~n861gat & ~n1068gat;
  assign n781 = n957gat & n861gat & ~n1068gat;
  assign n782 = ~n861gat & n1068gat & n957gat;
  assign n783 = ~n957gat & n861gat & n1068gat;
  assign n784_1 = ~n788 & ~n787 & ~n785 & ~n786;
  assign n785 = ~n1241gat & ~n1298gat & ~n1294gat;
  assign n786 = n1241gat & n1298gat & ~n1294gat;
  assign n787 = ~n1298gat & n1294gat & n1241gat;
  assign n788 = ~n1241gat & n1298gat & n1294gat;
  assign n789_1 = ~n784_1 & n774_1 & ~n779_1;
  assign n790 = ~n774_1 & n779_1 & ~n784_1;
  assign n791 = n784_1 & n774_1 & n779_1;
  assign n3120gat = n793 | n799_1;
  assign n793 = n716 & ~n794_1;
  assign n794_1 = ~n798 & ~n797 & ~n795 & ~n796;
  assign n795 = ~n584gat & n713;
  assign n796 = ~n865gat & n711;
  assign n797 = ~n322gat & n715;
  assign n798 = ~n341gat & n700;
  assign n799_1 = ~n818 & ~n817 & ~n800 & ~n816;
  assign n800 = n811 & ~n801 & ~n806;
  assign n801 = ~n805 & ~n804_1 & ~n802 & ~n803;
  assign n802 = ~n275gat & ~n398gat & ~n402gat;
  assign n803 = ~n275gat & n398gat & n402gat;
  assign n804_1 = ~n398gat & n402gat & n275gat;
  assign n805 = n275gat & n398gat & ~n402gat;
  assign n806 = ~n810 & ~n809_1 & ~n807 & ~n808;
  assign n807 = ~n165gat & ~n279gat & ~n283gat;
  assign n808 = n165gat & n279gat & ~n283gat;
  assign n809_1 = ~n279gat & n283gat & n165gat;
  assign n810 = ~n165gat & n279gat & n283gat;
  assign n811 = ~n815 & ~n814_1 & ~n812 & ~n813;
  assign n812 = ~n1026gat & ~n919gat & ~n846gat;
  assign n813 = n1026gat & n919gat & ~n846gat;
  assign n814_1 = ~n919gat & n846gat & n1026gat;
  assign n815 = ~n1026gat & n919gat & n846gat;
  assign n816 = ~n811 & n801 & ~n806;
  assign n817 = ~n801 & n806 & ~n811;
  assign n818 = n811 & n801 & n806;
  assign n3121gat = n820 | n826;
  assign n820 = n716 & ~n821;
  assign n821 = ~n825 & ~n824_1 & ~n822 & ~n823;
  assign n822 = ~n314gat & n715;
  assign n823 = ~n1148gat & n711;
  assign n824_1 = ~n699gat & n713;
  assign n825 = ~n394gat & n700;
  assign n826 = ~n845 & ~n844_1 & ~n827 & ~n843;
  assign n827 = n838 & ~n828 & ~n833;
  assign n828 = ~n832 & ~n831 & ~n829_1 & ~n830;
  assign n829_1 = ~n684gat & ~n699gat & ~n584gat;
  assign n830 = n684gat & n699gat & ~n584gat;
  assign n831 = ~n699gat & n584gat & n684gat;
  assign n832 = ~n684gat & n699gat & n584gat;
  assign n833 = ~n837 & ~n836 & ~n834_1 & ~n835;
  assign n834_1 = ~n816gat & ~n580gat & ~n680gat;
  assign n835 = n816gat & n580gat & ~n680gat;
  assign n836 = ~n580gat & n680gat & n816gat;
  assign n837 = ~n816gat & n580gat & n680gat;
  assign n838 = ~n842 & ~n841 & ~n839_1 & ~n840;
  assign n839_1 = ~n820gat & ~n883gat & ~n824gat;
  assign n840 = n820gat & n883gat & ~n824gat;
  assign n841 = ~n883gat & n824gat & n820gat;
  assign n842 = ~n820gat & n883gat & n824gat;
  assign n843 = ~n838 & n828 & ~n833;
  assign n844_1 = ~n828 & n833 & ~n838;
  assign n845 = n838 & n828 & n833;
  assign n3122gat = n847 | n853;
  assign n847 = n716 & ~n848;
  assign n848 = ~n852 & ~n851 & ~n849_1 & ~n850;
  assign n849_1 = ~n318gat & n715;
  assign n850 = ~n703gat & n700;
  assign n851 = ~n684gat & n713;
  assign n852 = ~n1080gat & n711;
  assign n853 = ~n872 & ~n871 & ~n854_1 & ~n870;
  assign n854_1 = n865 & ~n855 & ~n860;
  assign n855 = ~n859_1 & ~n858 & ~n856 & ~n857;
  assign n856 = ~n614gat & ~n491gat & ~n618gat;
  assign n857 = ~n614gat & n491gat & n618gat;
  assign n858 = ~n491gat & n618gat & n614gat;
  assign n859_1 = n614gat & n491gat & ~n618gat;
  assign n860 = ~n864_1 & ~n863 & ~n861 & ~n862;
  assign n861 = ~n707gat & ~n838gat & ~n834gat;
  assign n862 = n707gat & n838gat & ~n834gat;
  assign n863 = ~n838gat & n834gat & n707gat;
  assign n864_1 = ~n707gat & n838gat & n834gat;
  assign n865 = ~n869_1 & ~n868 & ~n866 & ~n867;
  assign n866 = ~n830gat & ~n626gat & ~n622gat;
  assign n867 = n830gat & n626gat & ~n622gat;
  assign n868 = ~n626gat & n622gat & n830gat;
  assign n869_1 = ~n830gat & n626gat & n622gat;
  assign n870 = ~n865 & n855 & ~n860;
  assign n871 = ~n855 & n860 & ~n865;
  assign n872 = n865 & n855 & n860;
  assign n3123gat = n874_1 | n880;
  assign n874_1 = n716 & ~n875;
  assign n875 = ~n879_1 & ~n878 & ~n876 & ~n877;
  assign n876 = ~n1294gat & n711;
  assign n877 = ~n726gat & n700;
  assign n878 = ~n561gat & n715;
  assign n879_1 = ~n824gat & n713;
  assign n880 = ~n881 & ~n900;
  assign n881 = ~n667gat & n882;
  assign n882 = ~n899_1 & ~n898 & ~n883 & ~n897;
  assign n883 = n894_1 & ~n884_1 & ~n889_1;
  assign n884_1 = ~n888 & ~n887 & ~n885 & ~n886;
  assign n885 = ~n318gat & ~n314gat & ~n322gat;
  assign n886 = n318gat & n314gat & ~n322gat;
  assign n887 = ~n314gat & n322gat & n318gat;
  assign n888 = ~n318gat & n314gat & n322gat;
  assign n889_1 = ~n893 & ~n892 & ~n890 & ~n891;
  assign n890 = ~n553gat & ~n777gat & ~n659gat;
  assign n891 = n553gat & n777gat & ~n659gat;
  assign n892 = ~n777gat & n659gat & n553gat;
  assign n893 = ~n553gat & n777gat & n659gat;
  assign n894_1 = ~n895 & ~n896;
  assign n895 = n561gat & ~n366gat;
  assign n896 = ~n561gat & n366gat;
  assign n897 = ~n894_1 & n884_1 & ~n889_1;
  assign n898 = ~n884_1 & n889_1 & ~n894_1;
  assign n899_1 = n894_1 & n884_1 & n889_1;
  assign n900 = n667gat & ~n882;
  assign n3124gat = n902 | n910;
  assign n902 = n716 & ~n903;
  assign n903 = ~n909_1 & ~n908 & ~n907 & ~n904_1 & ~n905;
  assign n904_1 = ~n883gat & n713;
  assign n905 = ~n673gat & n906;
  assign n906 = n704_1 & n707 & ~n701;
  assign n907 = ~n366gat & n715;
  assign n908 = ~n722gat & n700;
  assign n909_1 = ~n1298gat & n711;
  assign n910 = ~n911 & ~n912;
  assign n911 = n1197gat & ~n678;
  assign n912 = ~n1197gat & n678;
  assign n3125gat = n914_1 | n922;
  assign n914_1 = n716 & ~n915;
  assign n915 = ~n920 & ~n919_1 & ~n918 & ~n916 & ~n917 & ~n921;
  assign n916 = n715 & ~n882;
  assign n917 = ~n707 & n701 & n704_1;
  assign n918 = ~n1241gat & n711;
  assign n919_1 = n673gat & n906;
  assign n920 = ~n842gat & n700;
  assign n921 = ~n820gat & n713;
  assign n922 = ~n923 & ~n929_1;
  assign n923 = ~n926 & ~n924_1 & ~n925;
  assign n924_1 = n2495gat & n2390gat;
  assign n925 = ~n2495gat & ~n2390gat;
  assign n926 = ~n928 & ~n927 & ~n924_1 & ~n925;
  assign n927 = n2270gat & ~n2339gat;
  assign n928 = ~n2270gat & n2339gat;
  assign n929_1 = ~n926 & ~n927 & ~n928;
  assign n3129gat = n931 | n941;
  assign n931 = ~n915 & ~n932;
  assign n932 = ~n933 & ~n940;
  assign n933 = ~n934_1 & n935;
  assign n934_1 = n3088gat & n3093gat;
  assign n935 = ~n939_1 & ~n938 & ~n936 & ~n937;
  assign n936 = n934_1 & n708 & n702 & n705;
  assign n937 = ~n702 & ~n708;
  assign n938 = n3084gat & n3093gat;
  assign n939_1 = n3083gat & n3093gat;
  assign n940 = n709_1 & n703 & n717 & n706;
  assign n941 = ~n942 & ~n944_1;
  assign n942 = ~n716 & ~n943;
  assign n943 = n934_1 & n935;
  assign n944_1 = ~n947 & ~n945 & ~n946;
  assign n945 = ~n678 & n715;
  assign n946 = ~n830gat & n713;
  assign n947 = ~n1026gat & n711;
  assign n3130gat = n949_1 | n950;
  assign n949_1 = ~n698 & ~n932;
  assign n950 = ~n942 & ~n951;
  assign n951 = ~n954_1 & ~n952 & ~n953;
  assign n952 = ~n1035gat & n715;
  assign n953 = ~n283gat & n711;
  assign n954_1 = ~n834gat & n713;
  assign n3131gat = n956 | n961;
  assign n956 = ~n942 & ~n957;
  assign n957 = ~n960 & ~n958 & ~n959_1;
  assign n958 = ~n838gat & n713;
  assign n959_1 = ~n279gat & n711;
  assign n960 = ~n1072gat & n715;
  assign n961 = ~n740 & ~n932;
  assign n3132gat = n963 | n968;
  assign n963 = ~n942 & ~n964_1;
  assign n964_1 = ~n967 & ~n965 & ~n966;
  assign n965 = ~n707gat & n713;
  assign n966 = ~n165gat & n711;
  assign n967 = ~n1121gat & n715;
  assign n968 = ~n767 & ~n932;
  assign n3133gat = n970 | n971;
  assign n970 = ~n794_1 & ~n932;
  assign n971 = ~n942 & ~n972;
  assign n972 = ~n975 & ~n973 & ~n974_1;
  assign n973 = ~n614gat & n713;
  assign n974_1 = ~n275gat & n711;
  assign n975 = ~n931gat & n715;
  assign n3134gat = n977 | n982;
  assign n977 = ~n942 & ~n978;
  assign n978 = ~n981 & ~n979_1 & ~n980;
  assign n979_1 = ~n491gat & n713;
  assign n980 = ~n398gat & n711;
  assign n981 = ~n1045gat & n715;
  assign n982 = ~n821 & ~n932;
  assign n3135gat = n984_1 | n989_1;
  assign n984_1 = ~n942 & ~n985;
  assign n985 = ~n988 & ~n986 & ~n987;
  assign n986 = ~n1135gat & n715;
  assign n987 = ~n402gat & n711;
  assign n988 = ~n618gat & n713;
  assign n989_1 = ~n848 & ~n932;
  assign n3136gat = n991 | n992;
  assign n991 = ~n875 & ~n932;
  assign n992 = ~n942 & ~n993;
  assign n993 = ~n996 & ~n994_1 & ~n995;
  assign n994_1 = ~n622gat & n713;
  assign n995 = ~n846gat & n711;
  assign n996 = ~n1282gat & n715;
  assign n3137gat = n998 | n999_1;
  assign n998 = ~n903 & ~n932;
  assign n999_1 = ~n942 & ~n1000;
  assign n1000 = ~n1003 & ~n1001 & ~n1002;
  assign n1001 = ~n1226gat & n715;
  assign n1002 = ~n919gat & n711;
  assign n1003 = ~n626gat & n713;
  assign n3138gat = ~n1005 & n1009_1 & n1011;
  assign n1005 = ~n1006 & ~n1008;
  assign n1006 = n726gat & n722gat & n1007 & ~n2454gat;
  assign n1007 = n394gat & ~n703gat;
  assign n1008 = n726gat & ~n722gat & n1007 & ~n2454gat;
  assign n1009_1 = ~n2207gat & ~n2562gat & n1010 & ~n2203gat;
  assign n1010 = n2399gat & n2343gat;
  assign n1011 = n2543gat & n2490gat & ~n2626gat & n2622gat & n2630gat;
  assign n1012 = ~n1045 & ~n1043 & ~n1037 & ~n1013 & ~n1032 & ~n1046;
  assign n1013 = ~n1508gat & ~n1014_1;
  assign n1014_1 = ~n1015 & ~n1029_1;
  assign n1015 = ~n1016 & n1018;
  assign n1016 = ~n2203gat & n2399gat & n1017 & ~n2207gat;
  assign n1017 = ~n2343gat & n2562gat;
  assign n1018 = ~n1027 & ~n1019_1 & ~n1340gat;
  assign n1019_1 = n1020 & n1024_1;
  assign n1020 = ~n1021 & ~n1023;
  assign n1021 = n1022 & ~n722gat & ~n726gat;
  assign n1022 = ~n2454gat & n394gat & n703gat;
  assign n1023 = ~n726gat & n1022 & n722gat;
  assign n1024_1 = ~n1026 & n1005 & ~n1025;
  assign n1025 = ~n722gat & n726gat & n1022;
  assign n1026 = n703gat & ~n394gat & ~n2454gat & n722gat & n726gat;
  assign n1027 = n2102gat & ~n1028;
  assign n1028 = ~n1880gat & ~n1763gat;
  assign n1029_1 = ~n1462gat & n1030 & n1394gat;
  assign n1030 = ~n1027 & ~n1031;
  assign n1031 = n1767gat & n1880gat & n1834gat;
  assign n1032 = ~n1678gat & ~n1033;
  assign n1033 = ~n1034_1 & ~n1035;
  assign n1034_1 = n1462gat & ~n1027;
  assign n1035 = ~n1596gat & n1036;
  assign n1036 = ~n1020 & n1027;
  assign n1037 = n1871gat & ~n1775gat & ~n3098gat & ~n1038 & ~n1041;
  assign n1038 = n1825gat & ~n1039_1;
  assign n1039_1 = ~n1775gat & n1040 & n3097gat;
  assign n1040 = n1880gat & n2021gat;
  assign n1041 = ~n1829gat & n1042;
  assign n1042 = n1821gat & n1825gat;
  assign n1043 = ~n1525gat & n1044_1;
  assign n1044_1 = n1027 & ~n1024_1 & ~n1394gat;
  assign n1045 = ~n1596gat & n1394gat & ~n1678gat & n1020 & n1027;
  assign n1046 = ~n1588gat & n1027 & n1596gat;
  assign n1047 = ~n1055 & ~n1054 & ~n1048 & ~n1050;
  assign n1048 = ~n1456gat & ~n1049;
  assign n1049 = ~n1018 & ~n1030;
  assign n1050 = ~n1748gat & ~n1051;
  assign n1051 = ~n1053 & ~n1052 & ~n1036;
  assign n1052 = ~n1024_1 & n1336gat & n1027;
  assign n1053 = n1027 & ~n1031;
  assign n1054 = n1340gat & ~n1027 & ~n1807gat;
  assign n1055 = ~n1675gat & n1044_1;
  assign n3143gat = ~n1057 | n1139;
  assign n1057 = ~n1138 & ~n1137 & ~n1136 & ~n1058 & ~n1080;
  assign n1058 = ~n1020 & ~n1059;
  assign n1059 = ~n1071 & ~n1069 & ~n1068 & ~n1060 & ~n1065 & ~n1072 & ~n1074 & ~n1076 & ~n1078;
  assign n1060 = ~n1061 & n1064 & ~n2203gat & ~n2207gat;
  assign n1061 = ~n1062 & ~n1063;
  assign n1062 = n882 & n1021;
  assign n1063 = ~n882 & ~n1021;
  assign n1064 = n2562gat & n1010;
  assign n1065 = n1067 & n1066 & ~n322gat;
  assign n1066 = ~n2343gat & n2399gat & ~n2562gat;
  assign n1067 = n2203gat & ~n2207gat;
  assign n1068 = ~n2399gat & n1017 & ~n561gat & n1067;
  assign n1069 = n1067 & n1070 & ~n777gat;
  assign n1070 = ~n2562gat & n1010;
  assign n1071 = n1067 & n1064 & ~n659gat;
  assign n1072 = n1067 & n1073 & ~n553gat;
  assign n1073 = n2399gat & n1017;
  assign n1074 = n1067 & n1075 & ~n314gat;
  assign n1075 = ~n2399gat & n2343gat & n2562gat;
  assign n1076 = n1067 & n1077 & ~n318gat;
  assign n1077 = ~n2399gat & n2343gat & ~n2562gat;
  assign n1078 = n1067 & n1079 & ~n366gat;
  assign n1079 = ~n2562gat & ~n2343gat & ~n2399gat;
  assign n1080 = n1389gat & ~n1081;
  assign n1081 = ~n1099 & ~n1095 & ~n1091 & ~n1082 & ~n1087 & ~n1102 & ~n1106 & ~n1108 & ~n1112 & ~n1116 & ~n1120 & ~n1124 & ~n1128 & ~n1132;
  assign n1082 = ~n1083 & n1075 & n1086;
  assign n1083 = ~n1084 & ~n1085;
  assign n1084 = ~n707gat & n1031;
  assign n1085 = ~n165gat & ~n1031;
  assign n1086 = ~n2203gat & n2207gat;
  assign n1087 = ~n1088 & n1066 & n1086;
  assign n1088 = ~n1089 & ~n1090;
  assign n1089 = ~n838gat & n1031;
  assign n1090 = ~n279gat & ~n1031;
  assign n1091 = ~n1092 & n1073 & n1086;
  assign n1092 = ~n1093 & ~n1094;
  assign n1093 = ~n834gat & n1031;
  assign n1094 = ~n283gat & ~n1031;
  assign n1095 = ~n1096 & n1077 & n1086;
  assign n1096 = ~n1097 & ~n1098;
  assign n1097 = ~n614gat & n1031;
  assign n1098 = ~n275gat & ~n1031;
  assign n1099 = ~n1100 & n1070 & n1101;
  assign n1100 = n1020 & ~n1026;
  assign n1101 = n2203gat & n2207gat;
  assign n1102 = n1017 & ~n1103 & ~n2399gat & n1101;
  assign n1103 = ~n1104 & ~n1105;
  assign n1104 = ~n1148gat & ~n1031;
  assign n1105 = ~n699gat & n1031;
  assign n1106 = ~n1107 & n1064 & n1101;
  assign n1107 = n2084gat & ~n1026;
  assign n1108 = ~n1109 & n1079 & n1101;
  assign n1109 = ~n1110 & ~n1111;
  assign n1110 = ~n1080gat & ~n1031;
  assign n1111 = ~n684gat & n1031;
  assign n1112 = ~n1113 & n1070 & n1086;
  assign n1113 = ~n1114 & ~n1115;
  assign n1114 = ~n883gat & n1031;
  assign n1115 = ~n1298gat & ~n1031;
  assign n1116 = ~n1117 & n1064 & n1086;
  assign n1117 = ~n1118 & ~n1119;
  assign n1118 = ~n1294gat & ~n1031;
  assign n1119 = ~n824gat & n1031;
  assign n1120 = ~n1121 & n1075 & n1101;
  assign n1121 = ~n1122 & ~n1123;
  assign n1122 = ~n816gat & n1031;
  assign n1123 = ~n957gat & ~n1031;
  assign n1124 = ~n1125 & n1073 & n1101;
  assign n1125 = ~n1126 & ~n1127;
  assign n1126 = ~n1068gat & ~n1031;
  assign n1127 = ~n680gat & n1031;
  assign n1128 = ~n1129 & n1066 & n1101;
  assign n1129 = ~n1130 & ~n1131;
  assign n1130 = ~n580gat & n1031;
  assign n1131 = ~n861gat & ~n1031;
  assign n1132 = ~n1133 & n1077 & n1101;
  assign n1133 = ~n1134 & ~n1135;
  assign n1134 = ~n865gat & ~n1031;
  assign n1135 = ~n584gat & n1031;
  assign n1136 = ~n1678gat & n1053 & ~n1394gat;
  assign n1137 = n1871gat & ~n2592gat & ~n673gat;
  assign n1138 = ~n1508gat & n1030 & ~n1394gat;
  assign n1139 = ~n1140 & ~n1152;
  assign n1140 = n1141 & ~n1146;
  assign n1141 = ~n1145 & ~n1144 & ~n1142 & ~n1143;
  assign n1142 = ~n2490gat & n2626gat & ~n2622gat;
  assign n1143 = ~n2622gat & n2490gat & ~n2626gat;
  assign n1144 = n2622gat & ~n2490gat & ~n2626gat;
  assign n1145 = n2622gat & n2490gat & n2626gat;
  assign n1146 = n1141 & n1147;
  assign n1147 = ~n1151 & ~n1150 & ~n1148 & ~n1149;
  assign n1148 = ~n2634gat & ~n2543gat & ~n2630gat;
  assign n1149 = n2634gat & n2543gat & ~n2630gat;
  assign n1150 = ~n2543gat & n2630gat & n2634gat;
  assign n1151 = ~n2634gat & n2543gat & n2630gat;
  assign n1152 = n1147 & ~n1146;
  assign n3144gat = ~n1057 | n1154;
  assign n1154 = ~n1155 & ~n1167;
  assign n1155 = n1156 & ~n1161;
  assign n1156 = ~n1160 & ~n1159 & ~n1157 & ~n1158;
  assign n1157 = n2640gat & ~n2562gat & ~n2343gat;
  assign n1158 = ~n2640gat & n2562gat & ~n2343gat;
  assign n1159 = ~n2562gat & n2343gat & ~n2640gat;
  assign n1160 = n2640gat & n2562gat & n2343gat;
  assign n1161 = n1156 & n1162;
  assign n1162 = ~n1166 & ~n1165 & ~n1163 & ~n1164;
  assign n1163 = ~n2207gat & ~n2399gat & ~n2203gat;
  assign n1164 = n2399gat & n1067;
  assign n1165 = n2399gat & n1086;
  assign n1166 = ~n2399gat & n1101;
  assign n1167 = n1162 & ~n1161;
  assign n3145gat = n1019_1 & ~n1169;
  assign n1169 = n2514gat & n649_1;
  assign n3146gat = n2169gat & n2176gat & n2033gat & n2037gat & ~n1171 & n2095gat & n2110gat;
  assign n1171 = n2514gat & n649_1 & n1871gat;
  assign n1172 = n2450gat & n2446gat;
  assign n3150gat = n1174 | ~n1175;
  assign n1174 = ~n337gat & ~n2454gat;
  assign n1175 = ~n1176 & ~n1177;
  assign n1176 = ~n2061gat & ~n632;
  assign n1177 = n2061gat & n632;
  assign n3151gat = ~n1179 | n624_1 | n635;
  assign n1179 = ~n1180 & n2139gat & ~n1181;
  assign n1180 = n2139gat & ~n1899gat;
  assign n1181 = ~n2139gat & n1899gat;
  assign n1182 = ~n1183 & ~n1184;
  assign n1183 = n3072gat & n3093gat;
  assign n1184 = n3081gat & n3095gat;
  assign n245 = n703gat & n394gat & n722gat & n726gat;
  assign n255 = ~n3099gat & n2319gat;
  assign n299 = n1188 | n1189;
  assign n1188 = n3065gat & n3093gat;
  assign n1189 = n3074gat & n3095gat;
  assign n304 = n1191 | n1192;
  assign n1191 = n3076gat & n3095gat;
  assign n1192 = n3067gat & n3093gat;
  assign n309 = n1194 | n1195;
  assign n1194 = n3075gat & n3095gat;
  assign n1195 = n3066gat & n3093gat;
  assign n314 = n1197 | n1198;
  assign n1197 = n3071gat & n3093gat;
  assign n1198 = n3080gat & n3095gat;
  assign n319 = n1200 | n1201;
  assign n1200 = n3073gat & n3093gat;
  assign n1201 = n3082gat & n3095gat;
  assign n328 = n1203 | n1204;
  assign n1203 = n3068gat & n3093gat;
  assign n1204 = n3077gat & n3095gat;
  assign n333 = n1206 | n1207;
  assign n1206 = n3070gat & n3093gat;
  assign n1207 = n3079gat & n3095gat;
  assign n338 = n1209 | n1210;
  assign n1209 = n3069gat & n3093gat;
  assign n1210 = n3078gat & n3095gat;
  assign n364 = n1212 | n1221;
  assign n1212 = n1213 & ~n1216;
  assign n1213 = ~n1214 & ~n1215;
  assign n1214 = n628 & n641 & ~n627;
  assign n1215 = n3088gat & n3087gat & n647 & n636 & ~n638;
  assign n1216 = ~n1220 & ~n1217 & ~n1219;
  assign n1217 = ~n148gat & ~n1218;
  assign n1218 = n1008 & ~n156gat & ~n152gat;
  assign n1219 = n148gat & n1218 & ~n256gat;
  assign n1220 = n256gat & ~n148gat;
  assign n1221 = n3065gat & ~n1213;
  assign n369 = n1223 | n1224;
  assign n1223 = n3067gat & ~n1213;
  assign n1224 = n1213 & ~n1225;
  assign n1225 = ~n1228 & ~n1226 & ~n1227;
  assign n1226 = n152gat & n1008 & ~n156gat;
  assign n1227 = n156gat & ~n152gat;
  assign n1228 = ~n152gat & ~n1008;
  assign n374 = n1230 | n1234;
  assign n1230 = n1213 & ~n1231;
  assign n1231 = ~n1232 & ~n1233;
  assign n1232 = n256gat & n1218;
  assign n1233 = ~n256gat & ~n1218;
  assign n1234 = n3066gat & ~n1213;
  assign n379 = n1236 | n1243;
  assign n1236 = n1213 & ~n1237;
  assign n1237 = ~n1238 & ~n1242;
  assign n1238 = n470gat & ~n1239;
  assign n1239 = ~n1240 & ~n1241;
  assign n1240 = n1008 & n256gat & ~n152gat;
  assign n1241 = n156gat & n1008;
  assign n1242 = ~n470gat & n1239;
  assign n1243 = n3073gat & ~n1213;
  assign n384 = n1245 | n1248;
  assign n1245 = n1213 & ~n1246;
  assign n1246 = ~n1241 & ~n1247;
  assign n1247 = ~n156gat & ~n1008;
  assign n1248 = n3068gat & ~n1213;
  assign n394 = n1250 | n1252;
  assign n1250 = n3065gat & n1251;
  assign n1251 = ~n3088gat & n3087gat & n647 & n636 & ~n638;
  assign n1252 = n3074gat & n1214;
  assign n399 = n1254 | n1255;
  assign n1254 = n3067gat & n1251;
  assign n1255 = n3076gat & n1214;
  assign n404 = n1257 | n1258;
  assign n1257 = n3075gat & n1214;
  assign n1258 = n3066gat & n1251;
  assign n409 = n1267 | n1260 | n1266;
  assign n1260 = n1261 & ~n1262;
  assign n1261 = ~n1214 & ~n1251;
  assign n1262 = ~n1265 & ~n1263 & ~n1264;
  assign n1263 = ~n331gat & ~n1006;
  assign n1264 = ~n388gat & n1006 & n331gat;
  assign n1265 = ~n331gat & n388gat;
  assign n1266 = n3080gat & n1214;
  assign n1267 = n3071gat & n1251;
  assign n414 = n1277 | n1269 | n1276;
  assign n1269 = n1261 & ~n1270;
  assign n1270 = ~n1271 & ~n1275;
  assign n1271 = ~n463gat & n1272;
  assign n1272 = ~n1273 & ~n1274;
  assign n1273 = n327gat & n1006 & ~n331gat;
  assign n1274 = n388gat & n1006;
  assign n1275 = n463gat & ~n1272;
  assign n1276 = n3073gat & n1251;
  assign n1277 = n3082gat & n1214;
  assign n419 = n1283 | n1279 | n1282;
  assign n1279 = n1261 & ~n1280;
  assign n1280 = ~n1274 & ~n1281;
  assign n1281 = ~n388gat & ~n1006;
  assign n1282 = n3072gat & n1251;
  assign n1283 = n3081gat & n1214;
  assign n424 = n1285 | n1286;
  assign n1285 = n3077gat & n1214;
  assign n1286 = n3068gat & n1251;
  assign n429 = n1294 | n1288 | n1293;
  assign n1288 = n1261 & ~n1289;
  assign n1289 = ~n1290 & ~n1292;
  assign n1290 = n327gat & n1291;
  assign n1291 = ~n388gat & n1006 & ~n331gat;
  assign n1292 = ~n327gat & ~n1291;
  assign n1293 = n3070gat & n1251;
  assign n1294 = n3079gat & n1214;
  assign n434 = n1302 | n1296 | n1301;
  assign n1296 = n1261 & ~n1297;
  assign n1297 = ~n1300 & ~n1298 & ~n1299;
  assign n1298 = ~n384gat & ~n1291;
  assign n1299 = n384gat & n1291 & ~n327gat;
  assign n1300 = n327gat & ~n384gat;
  assign n1301 = n3069gat & n1251;
  assign n1302 = n3078gat & n1214;
  assign n444 = ~n662 & n459;
  assign n459 = n1305 & n634;
  assign n1305 = ~n1306 & ~n1309;
  assign n1306 = ~n1027 & n1307;
  assign n1307 = n668 & n1308;
  assign n1308 = ~n2407gat & n660;
  assign n1309 = n1308 & n1027 & n667;
  assign n634 = n2095gat & ~n1311 & ~n1314 & n2037gat;
  assign n1311 = ~n3100gat & ~n1312;
  assign n1312 = n2309gat & n1313;
  assign n1313 = n2506gat & n2502gat & n2588gat & n2510gat & n2658gat;
  assign n1314 = n2099gat & ~n1040;
  assign n449 = ~n666 & n459;
  assign n454 = ~n657 & n459;
  assign n464 = ~n651 & n459;
  assign n469 = n634 & n1319;
  assign n1319 = ~n1330 & ~n1328 & ~n1320 & ~n1325;
  assign n1320 = ~n1321 & n1322 & ~n1323 & ~n1324;
  assign n1321 = n1740gat & ~n1027;
  assign n1322 = n632 & ~n2061gat & n1850gat & n2143gat;
  assign n1323 = ~n2091gat & n1027 & ~n1496gat;
  assign n1324 = ~n1740gat & ~n1027;
  assign n1325 = n1323 & n1009;
  assign n1009 = ~n1899gat & ~n2061gat & n1327 & n2143gat;
  assign n1327 = n2139gat & n1850gat;
  assign n1328 = n1324 & n1329;
  assign n1329 = ~n1850gat & ~n1899gat & n2139gat & n2143gat & n2061gat;
  assign n1330 = n1321 & n1014;
  assign n1014 = ~n2061gat & n1850gat & ~n2143gat & n632;
  assign n474 = ~n1179 & n469;
  assign n479 = ~n1175 & n469;
  assign n484 = ~n629_1 & n469;
  assign n489 = ~n642 & n469;
  assign n494 = ~n271gat & ~n2454gat;
  assign n499 = n2117gat & ~n1338 & ~n2125gat;
  assign n1338 = ~n3100gat & ~n1172;
  assign n504 = n494 & n1340;
  assign n1340 = ~n1338 & n2472gat & ~n1041;
  assign n514 = n1342 | n1346;
  assign n1342 = n3065gat & ~n1343;
  assign n1343 = ~n1344 & ~n1345;
  assign n1344 = n641 & n627 & ~n628;
  assign n1345 = n3086gat & n3085gat & n637 & n636 & ~n638;
  assign n1346 = ~n1009_1 & ~n2207gat & ~n1016 & ~n1024_1 & ~n1347;
  assign n1347 = ~n1348 & ~n1349;
  assign n1348 = ~n2155gat & ~n2543gat & n2630gat & ~n2622gat & n2626gat & ~n2490gat;
  assign n1349 = n2155gat & n2630gat & ~n2622gat & ~n2626gat & n2490gat & n2543gat;
  assign n519 = n1346 | n1351;
  assign n1351 = n3067gat & ~n1343;
  assign n524 = n1346 | n1353;
  assign n1353 = n3066gat & ~n1343;
  assign n529 = n1346 | n1355;
  assign n1355 = n3071gat & ~n1343;
  assign n534 = n1346 | n1357;
  assign n1357 = n3072gat & ~n1343;
  assign n539 = n1346 | n1359;
  assign n1359 = n3068gat & ~n1343;
  assign n544 = n1346 | n1361;
  assign n1361 = n3070gat & ~n1343;
  assign n549 = n1346 | n1363;
  assign n1363 = n3069gat & ~n1343;
  assign n554 = n1346 | n1365;
  assign n1365 = n3073gat & ~n1343;
  assign n564 = n1369 | n1367 | n1346;
  assign n1367 = n3073gat & n1368;
  assign n1368 = n3093gat & ~n1346;
  assign n1369 = n3082gat & n1370;
  assign n1370 = n3095gat & ~n1346;
  assign n569 = n1373 | n1372 | n1346;
  assign n1372 = n3065gat & n1368;
  assign n1373 = n3074gat & n1370;
  assign n574 = n1376 | n1375 | n1346;
  assign n1375 = n3067gat & n1368;
  assign n1376 = n3076gat & n1370;
  assign n579 = n1379 | n1378 | n1346;
  assign n1378 = n3075gat & n1370;
  assign n1379 = n3066gat & n1368;
  assign n584 = n1382 | n1381 | n1346;
  assign n1381 = n3080gat & n1370;
  assign n1382 = n3071gat & n1368;
  assign n589 = n1385 | n1384 | n1346;
  assign n1384 = n3081gat & n1370;
  assign n1385 = n3072gat & n1368;
  assign n594 = n1388 | n1387 | n1346;
  assign n1387 = n3077gat & n1370;
  assign n1388 = n3068gat & n1368;
  assign n599 = n1391 | n1390 | n1346;
  assign n1390 = n3079gat & n1370;
  assign n1391 = n3070gat & n1368;
  assign n604 = n1394 | n1393 | n1346;
  assign n1393 = n3078gat & n1370;
  assign n1394 = n3069gat & n1368;
  assign n614 = ~n2599gat | ~n2464gat | ~n2522gat | n3090gat | ~n2518gat | ~n2476gat | ~n2468gat | ~n2526gat;
  assign n619 = n1400 | ~n459 | n1397;
  assign n1397 = ~n2644gat & n1398;
  assign n1398 = ~n1399 & ~n653 & ~n2440gat;
  assign n1399 = n2403gat & ~n2394gat;
  assign n1400 = n2644gat & ~n1398;
  assign n629 = n1403 | ~n634 | n1402;
  assign n1402 = n2266gat & ~n676;
  assign n1403 = ~n2266gat & n676;
  assign n639 = ~n675 & n634;
  assign n644 = ~n670 & n634;
  assign n654 = n1410 | ~n469 | n1407;
  assign n1407 = ~n1975gat & n1408;
  assign n1408 = ~n1409 & ~n631 & ~n1899gat;
  assign n1409 = n2061gat & ~n2139gat;
  assign n1410 = n1975gat & ~n1408;
  assign n664 = ~n726gat & ~n722gat & n1007 & ~n2454gat;
  assign n669 = ~n726gat & n722gat & n1007 & ~n2454gat;
  assign n729 = ~n1414 & n1417;
  assign n1414 = ~n1415 & ~n1416;
  assign n1415 = ~n1027 & n1329;
  assign n1416 = n1027 & n1322;
  assign n1417 = ~n2347gat & ~n2403gat & n668 & n2407gat;
  assign n734 = n669 | ~n1019_1 | n664;
  assign n739 = n2440gat & n2403gat & n2394gat & n2347gat & n1420 & ~n2407gat;
  assign n1420 = ~n1899gat & n2061gat & n1327 & n2143gat;
  assign n754 = n1850gat & ~n2139gat & ~n1899gat & n2061gat & n1417 & n2143gat;
  assign n784 = n1026 | ~n1020 | n1025;
  assign n789 = n1424 | n1425;
  assign n1424 = n672 & ~n1319 & ~n1305 & ~n2179gat & ~n2135gat;
  assign n1425 = ~n1305 & ~n1319 & ~n2182gat;
  assign n809 = n1340 & n669;
  assign n814 = ~n1447 & ~n1040 & n1428 & ~n1311;
  assign n1428 = ~n1441 & ~n1440 & ~n1439 & ~n1429 & ~n1437 & ~n1443 & ~n1444 & ~n1445 & ~n1446;
  assign n1429 = ~n1436 & n667 & n1435 & ~n1430 & n1433 & n1434;
  assign n1430 = ~n1431 & ~n1432;
  assign n1431 = ~n1031 & n1415;
  assign n1432 = n1053 & n1322;
  assign n1433 = n398gat & ~n919gat;
  assign n1434 = n398gat & ~n402gat;
  assign n1435 = n2347gat & ~n2407gat & ~n2403gat;
  assign n1436 = n398gat & ~n846gat;
  assign n1437 = ~n1430 & n1308 & n1438;
  assign n1438 = n2394gat & n2440gat;
  assign n1439 = n1434 & n668 & ~n1430 & n1436 & ~n1433 & n1435;
  assign n1440 = n1436 & n654_1 & n1435 & ~n1430 & n1433 & n1434;
  assign n1441 = ~n1434 & n1433 & n1436 & n1442 & ~n1430 & ~n2407gat & n654_1;
  assign n1442 = n2403gat & n2347gat;
  assign n1443 = ~n1434 & n668 & n1442 & ~n1430 & n1436 & ~n1433 & ~n2407gat;
  assign n1444 = n1438 & n1434 & ~n1430 & n1435 & ~n1436 & ~n1433;
  assign n1445 = ~n1434 & ~n1436 & n1438 & ~n1433 & ~n2407gat & ~n1430 & n1442 & n398gat;
  assign n1446 = n1442 & n667 & n1433 & ~n1430 & ~n2407gat & ~n1436 & ~n1434;
  assign n1447 = ~n1312gat & n1775gat;
  assign n824 = n1180 & ~n1027 & n644_1 & n1850gat;
  assign n829 = n1899gat & ~n2061gat & n1327 & n2143gat;
  assign n849 = n1451 | n1452;
  assign n1451 = n3086gat & n3085gat & ~n3088gat & n3087gat & n636 & ~n638;
  assign n1452 = n628 & n641 & n627;
  assign n864 = ~n2169gat & n1312gat & n1428 & ~n1311;
  assign n874 = ~n2040gat & ~n1316gat & ~n1775gat;
  assign n884 = ~n1040 & n1428;
  assign n994 = n1340 & n664;
  assign n999 = n2562gat & n2203gat & ~n2207gat & n1011 & n1010;
  assign n1004 = n1322 & n1428;
  assign n1019 = n1417 & n829;
  assign n1024 = n1415 & n1428 & ~n1307;
  assign n1029 = n1850gat & n2143gat & n1181 & n2061gat;
  assign n1034 = ~n2347gat & ~n2403gat & n2407gat & n1014 & n667;
  assign n1039 = ~n2347gat & ~n2403gat & n2407gat & n1322 & n667;
  assign n1044 = n1312gat & n1420;
  assign n3106gat = ~n1871gat;
  assign n3115gat = 1'b1;
  assign n3116gat = ~n678;
  assign n3126gat = ~n2339gat;
  assign n3127gat = ~n2270gat;
  assign n3128gat = ~n2390gat;
  assign n3139gat = ~n1012;
  assign n3140gat = ~n1012;
  assign n3141gat = ~n1047;
  assign n3142gat = ~n1047;
  assign n3147gat = ~n1172;
  assign n3148gat = ~n2450gat;
  assign n3149gat = ~n1031;
  assign n3152gat = 1'b1;
  assign n169 = ~n1182;
  assign n174 = n3069gat;
  assign n179 = n3070gat;
  assign n184 = n3072gat;
  assign n189 = n3071gat;
  assign n193 = n3069gat;
  assign n197 = n3070gat;
  assign n201 = n3072gat;
  assign n205 = n3071gat;
  assign n210 = ~n722;
  assign n215 = n3065gat;
  assign n220 = n3067gat;
  assign n225 = n3066gat;
  assign n230 = n3073gat;
  assign n235 = n3068gat;
  assign n240 = ~n745;
  assign n250 = ~n2472gat;
  assign n259 = n255;
  assign n264 = ~n1042;
  assign n269 = ~n2029gat;
  assign n273 = n3065gat;
  assign n277 = n3067gat;
  assign n281 = n3066gat;
  assign n285 = n3073gat;
  assign n289 = n3068gat;
  assign n294 = ~n799_1;
  assign n323 = ~n1182;
  assign n343 = ~n772;
  assign n347 = n3070gat;
  assign n351 = n3069gat;
  assign n355 = n3071gat;
  assign n359 = n3072gat;
  assign n389 = ~n853;
  assign n439 = ~n826;
  assign n509 = ~n1027;
  assign n559 = ~n910;
  assign n609 = ~n880;
  assign n624 = ~n1154;
  assign n649 = ~n922;
  assign n659 = ~n1139;
  assign n674 = ~n1031;
  assign n679 = ~n2543gat;
  assign n684 = ~n2622gat;
  assign n689 = ~n2490gat;
  assign n694 = ~n2626gat;
  assign n699 = ~n2630gat;
  assign n704 = ~n2399gat;
  assign n709 = ~n2343gat;
  assign n714 = ~n2562gat;
  assign n719 = ~n2207gat;
  assign n724 = ~n2203gat;
  assign n744 = ~n1394gat;
  assign n749 = ~n1024_1;
  assign n759 = ~n1332gat;
  assign n764 = ~n1005;
  assign n769 = ~n2270gat;
  assign n774 = ~n2339gat;
  assign n779 = ~n2390gat;
  assign n794 = ~n1433gat;
  assign n799 = ~n1316gat;
  assign n804 = ~n1363gat;
  assign n819 = ~n1775gat;
  assign n834 = 1'b1;
  assign n839 = ~n2309gat;
  assign n844 = ~n1313;
  assign n854 = ~n2095gat;
  assign n859 = ~n2176gat;
  assign n869 = ~n1019_1;
  assign n879 = ~n2044gat;
  assign n889 = ~n2025gat;
  assign n894 = ~n2495gat;
  assign n899 = ~n2037gat;
  assign n904 = ~n2033gat;
  assign n909 = ~n2110gat;
  assign n914 = ~n2125gat;
  assign n919 = ~n2121gat;
  assign n924 = ~n2634gat;
  assign n929 = ~n2640gat;
  assign n934 = ~n614gat;
  assign n939 = ~n707gat;
  assign n944 = ~n824gat;
  assign n949 = ~n883gat;
  assign n954 = ~n820gat;
  assign n959 = ~n684gat;
  assign n964 = ~n699gat;
  assign n969 = ~n838gat;
  assign n974 = ~n830gat;
  assign n979 = ~n834gat;
  assign n984 = ~n2592gat;
  assign n989 = ~n2458gat;
  always @ (posedge clock) begin
    n673gat <= n169;
    n398gat <= n174;
    n402gat <= n179;
    n919gat <= n184;
    n846gat <= n189;
    n394gat <= n193;
    n703gat <= n197;
    n722gat <= n201;
    n726gat <= n205;
    n2510gat <= n210;
    n271gat <= n215;
    n160gat <= n220;
    n337gat <= n225;
    n842gat <= n230;
    n341gat <= n235;
    n2522gat <= n240;
    n2472gat <= n245;
    n2319gat <= n250;
    n1821gat <= n255;
    n1825gat <= n259;
    n2029gat <= n264;
    n1829gat <= n269;
    n283gat <= n273;
    n165gat <= n277;
    n279gat <= n281;
    n1026gat <= n285;
    n275gat <= n289;
    n2476gat <= n294;
    n1068gat <= n299;
    n957gat <= n304;
    n861gat <= n309;
    n1294gat <= n314;
    n1241gat <= n319;
    n1298gat <= n323;
    n865gat <= n328;
    n1080gat <= n333;
    n1148gat <= n338;
    n2468gat <= n343;
    n618gat <= n347;
    n491gat <= n351;
    n622gat <= n355;
    n626gat <= n359;
    n834gat <= n364;
    n707gat <= n369;
    n838gat <= n374;
    n830gat <= n379;
    n614gat <= n384;
    n2526gat <= n389;
    n680gat <= n394;
    n816gat <= n399;
    n580gat <= n404;
    n824gat <= n409;
    n820gat <= n414;
    n883gat <= n419;
    n584gat <= n424;
    n684gat <= n429;
    n699gat <= n434;
    n2464gat <= n439;
    n2399gat <= n444;
    n2343gat <= n449;
    n2203gat <= n454;
    n2562gat <= n459;
    n2207gat <= n464;
    n2626gat <= n469;
    n2490gat <= n474;
    n2622gat <= n479;
    n2630gat <= n484;
    n2543gat <= n489;
    n2102gat <= n494;
    n1880gat <= n499;
    n1763gat <= n504;
    n2155gat <= n509;
    n1035gat <= n514;
    n1121gat <= n519;
    n1072gat <= n524;
    n1282gat <= n529;
    n1226gat <= n534;
    n931gat <= n539;
    n1135gat <= n544;
    n1045gat <= n549;
    n1197gat <= n554;
    n2518gat <= n559;
    n667gat <= n564;
    n659gat <= n569;
    n553gat <= n574;
    n777gat <= n579;
    n561gat <= n584;
    n366gat <= n589;
    n322gat <= n594;
    n318gat <= n599;
    n314gat <= n604;
    n2599gat <= n609;
    n2588gat <= n614;
    n2640gat <= n619;
    n2658gat <= n624;
    n2495gat <= n629;
    n2390gat <= n634;
    n2270gat <= n639;
    n2339gat <= n644;
    n2502gat <= n649;
    n2634gat <= n654;
    n2506gat <= n659;
    n1834gat <= n664;
    n1767gat <= n669;
    n2084gat <= n674;
    n2143gat <= n679;
    n2061gat <= n684;
    n2139gat <= n689;
    n1899gat <= n694;
    n1850gat <= n699;
    n2403gat <= n704;
    n2394gat <= n709;
    n2440gat <= n714;
    n2407gat <= n719;
    n2347gat <= n724;
    n1389gat <= n729;
    n2021gat <= n734;
    n1394gat <= n739;
    n1496gat <= n744;
    n2091gat <= n749;
    n1332gat <= n754;
    n1740gat <= n759;
    n2179gat <= n764;
    n2190gat <= n769;
    n2135gat <= n774;
    n2262gat <= n779;
    n2182gat <= n784;
    n1433gat <= n789;
    n1316gat <= n794;
    n1363gat <= n799;
    n1312gat <= n804;
    n1775gat <= n809;
    n1871gat <= n814;
    n2592gat <= n819;
    n1508gat <= n824;
    n1678gat <= n829;
    n2309gat <= n834;
    n2450gat <= n839;
    n2446gat <= n844;
    n2095gat <= n849;
    n2176gat <= n854;
    n2169gat <= n859;
    n2454gat <= n864;
    n2040gat <= n869;
    n2044gat <= n874;
    n2037gat <= n879;
    n2025gat <= n884;
    n2099gat <= n889;
    n2266gat <= n894;
    n2033gat <= n899;
    n2110gat <= n904;
    n2125gat <= n909;
    n2121gat <= n914;
    n2117gat <= n919;
    n1975gat <= n924;
    n2644gat <= n929;
    n156gat <= n934;
    n152gat <= n939;
    n331gat <= n944;
    n388gat <= n949;
    n463gat <= n954;
    n327gat <= n959;
    n384gat <= n964;
    n256gat <= n969;
    n470gat <= n974;
    n148gat <= n979;
    n2458gat <= n984;
    n2514gat <= n989;
    n1771gat <= n994;
    n1336gat <= n999;
    n1748gat <= n1004;
    n1675gat <= n1009;
    n1807gat <= n1014;
    n1340gat <= n1019;
    n1456gat <= n1024;
    n1525gat <= n1029;
    n1462gat <= n1034;
    n1596gat <= n1039;
    n1588gat <= n1044;
  end
endmodule


