module medium_3 ( clock, 
    g43, g49, g633, g634, g635, g645, g647, g648, g690, g694, g698, g702,
    g722, g723, g751, g752, g753, g754, g755, g756, g757, g781, g941, g962,
    g1000, g1008, g1016, g1080, g1234, g1553, g1554, g786, g1206, g929,
    g955, g795, g1194, g1198, g1202, g24, g1203, g1196, g29, g22, g28, g10,
    g23, g37, g26, g1, g27, g42, g11, g32, g41, g31, g45, g9, g44, g21,
    g30, g25,
    g206, g291, g372, g453, g534, g594, g785, g1006, g1015, g1017, g1246,
    g1724, g1783, g1798, g1804, g1810, g1817, g1824, g1829, g1870, g1871,
    g1894, g1911, g1944, g2662, g2844, g2888, g3077, g3096, g3130, g3159,
    g3191, g3829, g3859, g3860, g4267, g4316, g4370, g4371, g4372, g4373,
    g4655, g4657, g4660, g4661, g4663, g4664, g5143, g5164, g5571, g5669,
    g5678, g5682, g5684, g5687, g5729, g6207, g6212, g6223, g6236, g6269,
    g6425, g6648, g6653, g6675, g6849, g6850, g6895, g6909, g7048, g7063,
    g7103, g7283, g7284, g7285, g7286, g7287, g7288, g7289, g7290, g7291,
    g7292, g7293, g7294, g7295, g7298, g7423, g7424, g7425, g7474, g7504,
    g7505, g7506, g7507, g7508, g7514, g7729, g7730, g7731, g7732, g8216,
    g8217, g8218, g8219, g8234, g8661, g8663, g8872, g8958, g9128, g9132,
    g9204, g9280, g9297, g9299, g9305, g9308, g9310, g9312, g9314, g9378,
    g7763, g1205, g3856, g3857, g3854, g1193, g1197, g1201, g6294, g6376,
    g1195, g6300, g6292, g6298, g6291, g6293, g6304, g6296, g6289, g6297,
    g6306, g6290, g6303, g6305, g6302, g6308, g6288, g6307, g6299, g6301,
    g6295  );
  input  clock, g43, g49, g633, g634, g635, g645, g647, g648, g690, g694, g698,
    g702, g722, g723, g751, g752, g753, g754, g755, g756, g757, g781, g941,
    g962, g1000, g1008, g1016, g1080, g1234, g1553, g1554, g786, g1206,
    g929, g955, g795, g1194, g1198, g1202, g24, g1203, g1196, g29, g22,
    g28, g10, g23, g37, g26, g1, g27, g42, g11, g32, g41, g31, g45, g9,
    g44, g21, g30, g25;
  output g206, g291, g372, g453, g534, g594, g785, g1006, g1015, g1017, g1246,
    g1724, g1783, g1798, g1804, g1810, g1817, g1824, g1829, g1870, g1871,
    g1894, g1911, g1944, g2662, g2844, g2888, g3077, g3096, g3130, g3159,
    g3191, g3829, g3859, g3860, g4267, g4316, g4370, g4371, g4372, g4373,
    g4655, g4657, g4660, g4661, g4663, g4664, g5143, g5164, g5571, g5669,
    g5678, g5682, g5684, g5687, g5729, g6207, g6212, g6223, g6236, g6269,
    g6425, g6648, g6653, g6675, g6849, g6850, g6895, g6909, g7048, g7063,
    g7103, g7283, g7284, g7285, g7286, g7287, g7288, g7289, g7290, g7291,
    g7292, g7293, g7294, g7295, g7298, g7423, g7424, g7425, g7474, g7504,
    g7505, g7506, g7507, g7508, g7514, g7729, g7730, g7731, g7732, g8216,
    g8217, g8218, g8219, g8234, g8661, g8663, g8872, g8958, g9128, g9132,
    g9204, g9280, g9297, g9299, g9305, g9308, g9310, g9312, g9314, g9378,
    g7763, g1205, g3856, g3857, g3854, g1193, g1197, g1201, g6294, g6376,
    g1195, g6300, g6292, g6298, g6291, g6293, g6304, g6296, g6289, g6297,
    g6306, g6290, g6303, g6305, g6302, g6308, g6288, g6307, g6299, g6301,
    g6295;
  reg g397, g1271, g312, g273, g452, g948, g629, g207, g1541, g1153, g940,
    g976, g498, g314, g1092, g454, g196, g535, g292, g772, g1375, g689,
    g183, g359, g1384, g1339, g20, g1424, g767, g393, g1077, g1231, g294,
    g1477, g4, g608, g1205, g465, g774, g921, g1304, g243, g1499, g80,
    g1444, g1269, g600, g423, g771, g803, g843, g315, g455, g906, g622,
    g891, g1014, g984, g117, g137, g527, g1513, g278, g1378, g718, g598,
    g1182, g1288, g1382, g179, g624, g48, g362, g878, g270, g763, g710,
    g730, g295, g1037, g1102, g483, g775, g621, g1364, g1454, g1296, g5,
    g1532, g587, g741, g13, g606, g1012, g52, g646, g1412, g327, g1189,
    g1389, g1029, g1371, g1429, g398, g985, g354, g619, g113, g133, g180,
    g1138, g1309, g889, g390, g625, g417, g681, g437, g351, g1201, g109,
    g1049, g1098, g200, g240, g479, g126, g596, g1268, g222, g420, g3, g58,
    g172, g387, g840, g365, g1486, g1504, g1185, g1385, g583, g822, g1025,
    g969, g768, g174, g685, g1087, g355, g911, g1226, g99, g1045, g1173,
    g1373, g186, g760, g959, g1369, g1007, g1459, g758, g480, g396, g612,
    g38, g632, g1415, g1227, g246, g449, g517, g118, g138, g16, g284, g142,
    g219, g426, g1388, g806, g846, g1428, g579, g1030, g614, g1430, g1247,
    g669, g110, g130, g225, g281, g819, g1308, g611, g631, g1217, g104,
    g1365, g825, g1333, g474, g1396, g141, g1509, g766, g1018, g588, g1467,
    g317, g457, g486, g471, g1381, g1197, g513, g1397, g533, g1021, g1421,
    g952, g1263, g580, g615, g1257, g46, g402, g998, g1041, g297, g954,
    g105, g145, g212, g1368, g232, g990, g475, g33, g951, g799, g812, g567,
    g313, g333, g168, g214, g234, g652, g1126, g1400, g1326, g92, g309,
    g211, g834, g231, g557, g1383, g1220, g158, g627, g661, g77, g831,
    g1327, g293, g1146, g89, g150, g773, g859, g1240, g518, g1472, g1443,
    g436, g405, g1034, g1147, g374, g98, g563, g510, g530, g215, g235,
    g1013, g6, g55, g1317, g504, g665, g544, g371, g62, g792, g468, g815,
    g1460, g553, g623, g501, g1190, g1390, g74, g1156, g318, g458, g342,
    g1250, g1163, g1363, g1432, g1053, g252, g330, g264, g1157, g1357,
    g375, g68, g852, g261, g516, g536, g979, g778, g199, g1292, g290,
    g1084, g1439, g770, g1276, g890, g1004, g1404, g93, g2, g287, g560,
    g1224, g1320, g617, g316, g336, g933, g456, g345, g628, g8, g887, g789,
    g173, g550, g255, g949, g1244, g620, g1435, g477, g926, g368, g855,
    g1214, g1110, g1310, g296, g972, g1402, g1236, g896, g613, g566, g1394,
    g1489, g883, g47, g971, g609, g103, g1254, g556, g1409, g626, g1229,
    g782, g237, g942, g228, g706, g746, g1462, g963, g129, g837, g599,
    g1192, g828, g1392, g492, g95, g944, g195, g1431, g1252, g356, g953,
    g1176, g1376, g1005, g1405, g901, g1270, g1225, g1073, g1324, g1069,
    g443, g1377, g377, g618, g602, g213, g233, g1199, g1399, g83, g888,
    g573, g399, g1245, g507, g547, g108, g610, g630, g1207, g249, g65,
    g916, g936, g478, g604, g945, g1114, g100, g429, g809, g849, g1408,
    g1336, g601, g122, g1065, g1122, g1228, g495, g1322, g1230, g1033,
    g267, g1195, g1395, g373, g274, g1266, g714, g734, g1142, g1342, g769,
    g1081, g1481, g1097, g543, g1154, g1354, g489, g874, g121, g591, g616,
    g1267, g1312, g605, g182, g1401, g950, g1329, g408, g871, g759, g146,
    g202, g440, g476, g184, g1149, g1398, g210, g394, g86, g570, g275,
    g303, g125, g181, g1524, g595, g1319, g863, g1211, g966, g1186, g1386,
    g875, g1170, g1370, g201, g1325, g1280, g1106, g1061, g1387, g762,
    g1461, g378, g1200, g1514, g1403, g1345, g1191, g1391, g185, g1307,
    g1159, g1223, g446, g1416, g395, g764, g1251, g216, g236, g205, g540,
    g576, g1537, g727, g999, g761, g1272, g1243, g1328, g1130, g1330, g114,
    g134, g1166, g524, g1366, g348, g1148, g1348, g1155, g1260, g7, g258,
    g521, g300, g765, g1118, g1167, g1318, g1367, g677, g376, g1057, g973,
    g1193, g1393, g1549, g1321, g1253, g1519, g584, g539, g324, g432,
    g1158, g321, g1311, g414, g1374, g94, g1284, g1545, g1380, g673, g607,
    g306, g943, g162, g411, g866, g1204, g1300, g384, g339, g459, g1323,
    g381, g1528, g1351, g597, g1372, g154, g435, g970, g1134, g995, g190,
    g1313, g603, g1494, g462, g1160, g1360, g1450, g187, g1179, g1379, g12,
    g71;
  wire n2131, n2132, n2139, n2141, n2142, n2151, n2152, n2153, n2154,
    n2155_1, n2156, n2157, n2158, n2159, n2160_1, n2161, n2162, n2163,
    n2164, n2165_1, n2166, n2167, n2168, n2169, n2170_1, n2171, n2172,
    n2173, n2174, n2175_1, n2179, n2180_1, n2181, n2190_1, n2191, n2196,
    n2200_1, n2201, n2202, n2203, n2205_1, n2206, n2208, n2209, n2212,
    n2213, n2214, n2215_1, n2216, n2217, n2219, n2220_1, n2221, n2222,
    n2223, n2224, n2225_1, n2226, n2227, n2228, n2229_1, n2230, n2231,
    n2232, n2233, n2234_1, n2235, n2236, n2237, n2238_1, n2239, n2240,
    n2241, n2242, n2243_1, n2244, n2245, n2246, n2247, n2248_1, n2249,
    n2250, n2251, n2252_1, n2253, n2254, n2255, n2256, n2257_1, n2258,
    n2259, n2260, n2261, n2262_1, n2263, n2264, n2265, n2266, n2267_1,
    n2268, n2269, n2270, n2271_1, n2272, n2273, n2274_1, n2275, n2276,
    n2277, n2278, n2279_1, n2280, n2281, n2282, n2283, n2284_1, n2285,
    n2286, n2287, n2288, n2289_1, n2290, n2291, n2292, n2293, n2294_1,
    n2295, n2296, n2297, n2298_1, n2299, n2300, n2301, n2302, n2303_1,
    n2304, n2305, n2306, n2307, n2308_1, n2309, n2310, n2311, n2312,
    n2313_1, n2314, n2315, n2316, n2317, n2318_1, n2319, n2322, n2323_1,
    n2324, n2325, n2326, n2327, n2328_1, n2329, n2330, n2331, n2332,
    n2333_1, n2334, n2335, n2336, n2337, n2338_1, n2339, n2340, n2341,
    n2342, n2343_1, n2344, n2345, n2346, n2347, n2348_1, n2349, n2350,
    n2351, n2352, n2353_1, n2354, n2355, n2356, n2357, n2358_1, n2359,
    n2360, n2361, n2364, n2365, n2366, n2367, n2368_1, n2369, n2370, n2371,
    n2372, n2373_1, n2374, n2375, n2376, n2377, n2378_1, n2379, n2380,
    n2381, n2382, n2383_1, n2384, n2385, n2386, n2387, n2388_1, n2389,
    n2390, n2391, n2392, n2393_1, n2394, n2395, n2396, n2397, n2398_1,
    n2399, n2400, n2401, n2402, n2405, n2406, n2407, n2408_1, n2409, n2410,
    n2411, n2412, n2413_1, n2414, n2415, n2416, n2417, n2418_1, n2419,
    n2420, n2421, n2422, n2423_1, n2424, n2425, n2426, n2427, n2428_1,
    n2429, n2430, n2431, n2432, n2433_1, n2434, n2435, n2436, n2437,
    n2438_1, n2439, n2440, n2441, n2444, n2445, n2446, n2447, n2448_1,
    n2449, n2450, n2451, n2452, n2453_1, n2454, n2455, n2456, n2457,
    n2458_1, n2459, n2460, n2461, n2462, n2463_1, n2464, n2465, n2466,
    n2467_1, n2468, n2469, n2470, n2471_1, n2472, n2473, n2474, n2475_1,
    n2476, n2477, n2478_1, n2479, n2480, n2483, n2484, n2485, n2486,
    n2487_1, n2488, n2489, n2490, n2491, n2492_1, n2493, n2494, n2495,
    n2496, n2497_1, n2498, n2499, n2500, n2501, n2502_1, n2503, n2504,
    n2505, n2506, n2507_1, n2508, n2509, n2510, n2513, n2514, n2515, n2516,
    n2517_1, n2518, n2519, n2520, n2521, n2522_1, n2523, n2524, n2525,
    n2526, n2527_1, n2528, n2529, n2530, n2531, n2532_1, n2533, n2534,
    n2535, n2536, n2537_1, n2538, n2539, n2540, n2543, n2544, n2545, n2546,
    n2547_1, n2548, n2549, n2550, n2551, n2552_1, n2553, n2554, n2555,
    n2556, n2557_1, n2558, n2559, n2560, n2561, n2562_1, n2563, n2564,
    n2565, n2566_1, n2567, n2568, n2569, n2572, n2574, n2575, n2576_1,
    n2577, n2578, n2579, n2580, n2581_1, n2582, n2583, n2584, n2585,
    n2586_1, n2587, n2588, n2589, n2590, n2591_1, n2592, n2593, n2594,
    n2595, n2596_1, n2597, n2598, n2599, n2600, n2601_1, n2602, n2603,
    n2604, n2605, n2606_1, n2607, n2608, n2609, n2610_1, n2611, n2612,
    n2613, n2614_1, n2615, n2616, n2617, n2618, n2620, n2621, n2622, n2623,
    n2624_1, n2625, n2629_1, n2630, n2631, n2632, n2634_1, n2635, n2636,
    n2637, n2638_1, n2639, n2641, n2642, n2644, n2645, n2648_1, n2649,
    n2651, n2652, n2653_1, n2654, n2655, n2657, n2658_1, n2659, n2660,
    n2662, n2663_1, n2665, n2666, n2667, n2668_1, n2669, n2670, n2671,
    n2672, n2673_1, n2674, n2675, n2676, n2677, n2679, n2680, n2681,
    n2683_1, n2684, n2686, n2687, n2688_1, n2689, n2690, n2691, n2693_1,
    n2694, n2695, n2696, n2697, n2698_1, n2699, n2700, n2701, n2702,
    n2703_1, n2704, n2705, n2706, n2707, n2708_1, n2709, n2710, n2711,
    n2712, n2713_1, n2714, n2715, n2716, n2717, n2718_1, n2719, n2720,
    n2721, n2722_1, n2723, n2724, n2725, n2729, n2730, n2731, n2732_1,
    n2733, n2734, n2735, n2736, n2737_1, n2738, n2739, n2740, n2741, n2743,
    n2744, n2745, n2747_1, n2748, n2749, n2751, n2752_1, n2753, n2755,
    n2756, n2758, n2760, n2761, n2763, n2764, n2765, n2766, n2767_1, n2768,
    n2769, n2770, n2771_1, n2774, n2775_1, n2777, n2778, n2780_1, n2781,
    n2783, n2784_1, n2785, n2787, n2788, n2789_1, n2791, n2792, n2793,
    n2794_1, n2795, n2796, n2798, n2799_1, n2801, n2802, n2804_1, n2805,
    n2807, n2808, n2810, n2811, n2813, n2814_1, n2815, n2817, n2818,
    n2819_1, n2821, n2822, n2824_1, n2826, n2827, n2829, n2830, n2831,
    n2832, n2833_1, n2835, n2836, n2837_1, n2838, n2840, n2841, n2842_1,
    n2844, n2845, n2846, n2847_1, n2848, n2850, n2851, n2852_1, n2853,
    n2855, n2857_1, n2858, n2860, n2861, n2862_1, n2863, n2864, n2865,
    n2866, n2867_1, n2868, n2869, n2870, n2871, n2872_1, n2873, n2874,
    n2875, n2876, n2877_1, n2878, n2879, n2880, n2881, n2882_1, n2883,
    n2886, n2887_1, n2889, n2890, n2891, n2892_1, n2893, n2895, n2896_1,
    n2897, n2899, n2900, n2901_1, n2903, n2904, n2905, n2906_1, n2907,
    n2908, n2909, n2910, n2912, n2913, n2914, n2916_1, n2917, n2919, n2920,
    n2921_1, n2923, n2924, n2926_1, n2927, n2929, n2930, n2931_1, n2933,
    n2934, n2936_1, n2937, n2940, n2941_1, n2943, n2944, n2946, n2947,
    n2949, n2950_1, n2952, n2953, n2954, n2955_1, n2957, n2958, n2960_1,
    n2961, n2963, n2964, n2966, n2967, n2968_1, n2969, n2970, n2972,
    n2973_1, n2974, n2976, n2977, n2979, n2981, n2982_1, n2983, n2984,
    n2985, n2986, n2988, n2989, n2991_1, n2992, n2994, n2995, n2997, n2998,
    n3000, n3002, n3003, n3005, n3006_1, n3007, n3008, n3009, n3012, n3013,
    n3014, n3015, n3017, n3018, n3020, n3021_1, n3023, n3024, n3026_1,
    n3027, n3029, n3030, n3032, n3033, n3036, n3038, n3039_1, n3041, n3042,
    n3044, n3045, n3047_1, n3048, n3049, n3052_1, n3053, n3054, n3055_1,
    n3057, n3058, n3060_1, n3061, n3063, n3065_1, n3066, n3068, n3069_1,
    n3070, n3072, n3073, n3075, n3076, n3077, n3079_1, n3080, n3082, n3083,
    n3085, n3086, n3088, n3089_1, n3091, n3092, n3093, n3096, n3097,
    n3099_1, n3100, n3102, n3103, n3104_1, n3106, n3108, n3109_1, n3111,
    n3113, n3114_1, n3116, n3117, n3119_1, n3120, n3122, n3124_1, n3126,
    n3127, n3130, n3131, n3132, n3134, n3135, n3137, n3138_1, n3140, n3141,
    n3143_1, n3144, n3145, n3146, n3148_1, n3149, n3150, n3151, n3152,
    n3153_1, n3154, n3156, n3157, n3159, n3160, n3162, n3163_1, n3165,
    n3166, n3167, n3168_1, n3169, n3171, n3172, n3174, n3175, n3177,
    n3178_1, n3179, n3180, n3181, n3182, n3183_1, n3185, n3186, n3188_1,
    n3189, n3190, n3192, n3193_1, n3195, n3197, n3198_1, n3200, n3201,
    n3202_1, n3204, n3205, n3207_1, n3208, n3210, n3211_1, n3212, n3213,
    n3215_1, n3216, n3218, n3219, n3221, n3222, n3224, n3225_1, n3226,
    n3228, n3229, n3232, n3234, n3235_1, n3237, n3238, n3240_1, n3241,
    n3242, n3243, n3244, n3245_1, n3246, n3247, n3248, n3250, n3251,
    n3253_1, n3254, n3257, n3258_1, n3260, n3261, n3263_1, n3264, n3265,
    n3266, n3267, n3268_1, n3270, n3271, n3273_1, n3274, n3276, n3277,
    n3279, n3280, n3282_1, n3283, n3284, n3285, n3286_1, n3288, n3289,
    n3291, n3292, n3294, n3295_1, n3297, n3298, n3299, n3301, n3302, n3303,
    n3304, n3306, n3308, n3309, n3310_1, n3312, n3313, n3316, n3317, n3319,
    n3320_1, n3321, n3322, n3324, n3325_1, n3326, n3327, n3328, n3329_1,
    n3330, n3332, n3333, n3335, n3336, n3338_1, n3339, n3341, n3342_1,
    n3343, n3344, n3345, n3346, n3347_1, n3348, n3350, n3351, n3353, n3354,
    n3356_1, n3357, n3359, n3360, n3362, n3363, n3366_1, n3367, n3369,
    n3370, n3372, n3373, n3374, n3375, n3377, n3378, n3379, n3380, n3381_1,
    n3382, n3383, n3384, n3385, n3386_1, n3387, n3388, n3389, n3390,
    n3391_1, n3392, n3393, n3394, n3395, n3396_1, n3397, n3398, n3399,
    n3400, n3401_1, n3402, n3403, n3405_1, n3406, n3407, n3410, n3411,
    n3413, n3414_1, n3415, n3416, n3417, n3418, n3420, n3421, n3423,
    n3424_1, n3426, n3427, n3429_1, n3430, n3432, n3433, n3434_1, n3435,
    n3437, n3438, n3440, n3441, n3443, n3444_1, n3446, n3448, n3449_1,
    n3451, n3452, n3455, n3456, n3458, n3460, n3461, n3462, n3463, n3465,
    n3466, n3468_1, n3469, n3470, n3471, n3472, n3473_1, n3474, n3476,
    n3477, n3478_1, n3480, n3481, n3483, n3484, n3486, n3487_1, n3489,
    n3490, n3492_1, n3493, n3495, n3496, n3498, n3499, n3502_1, n3503,
    n3507, n3508, n3510_1, n3511, n3512, n3514, n3515_1, n3517, n3518,
    n3521, n3523, n3524_1, n3526, n3527, n3528, n3530, n3531, n3532, n3533,
    n3535, n3536, n3538, n3539_1, n3540, n3541, n3542, n3543, n3544, n3546,
    n3547, n3548, n3549, n3550, n3551, n3553, n3554, n3556, n3557, n3560,
    n3561, n3563, n3564, n3566, n3567, n3569, n3571, n3572, n3574, n3576,
    n3578, n3579, n3581, n3582, n3585, n3586, n3588, n3589, n3591, n3592,
    n3594, n3595, n3597, n3598, n3599, n3600, n3602, n3603, n3605, n3607,
    n3608, n3610, n3611, n3613, n3614, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3624, n3625, n3626, n3629, n3630, n3633, n3634, n3636,
    n3637, n3638, n3639, n3640, n3641, n3642, n3644, n3645, n3647, n3648,
    n3650, n3651, n3653, n3654, n3657, n3658, n3660, n3661, n3663, n3664,
    n3666, n3667, n3668, n3669, n3671, n3672, n3674, n3676, n3677, n3679,
    n3680, n3682, n3683, n3685, n3686, n3689, n3691, n3692, n3693, n3694,
    n3695, n3696, n3697, n3699, n3700, n3701, n3704, n3705, n3707, n3708,
    n3710, n3711, n3713, n3714, n3715, n3718, n3719, n3721, n3722, n3724,
    n3725, n3727, n3728, n3730, n3731, n3732, n3733, n3735, n3736, n3738,
    n3739, n3741, n3744, n3745, n3747, n3748, n3749, n3750, n3751, n3752,
    n3753, n3755, n3757, n3758, n3760, n3761, n3763, n3764, n3766, n3767,
    n3769, n3770, n3772, n3773, n3775, n3776, n3777, n3778, n3779, n3781,
    n3782, n3784, n3785, n3787, n3788, n3790, n3791, n3793, n3794, n3796,
    n3797, n3799, n3800, n3803, n3804, n3805, n3807, n3808, n3810, n3811,
    n3813, n3814, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3824,
    n3825, n3827, n3828, n3830, n3831, n3832, n3833, n3834, n3836, n3837,
    n3839, n3840, n3841, n3843, n3845, n3846, n3848, n3849, n3851, n3853,
    n3854, n3856, n3857, n3859, n3860, n3862, n3863, n3864, n3865, n3867,
    n3868, n430, n435, n440, n445, n450, n455, n460, n465, n470, n475,
    n480, n485, n490, n495, n500, n505, n510, n515, n520, n525, n530, n535,
    n540, n545, n550, n555, n560, n565, n570, n575, n580, n585, n590, n595,
    n600, n605, n610, n614, n619, n624, n629, n634, n639, n644, n649, n654,
    n659, n664, n669, n674, n679, n684, n689, n694, n699, n704, n709, n714,
    n719, n724, n729, n734, n739, n744, n749, n754, n759, n764, n769, n774,
    n779, n784, n789, n794, n799, n804, n809, n814, n819, n824, n829, n834,
    n839, n844, n849, n854, n859, n864, n869, n874, n879, n884, n889, n894,
    n898, n903, n908, n913, n918, n923, n928, n933, n938, n943, n948, n953,
    n958, n963, n968, n973, n978, n983, n988, n993, n998, n1003, n1008,
    n1013, n1018, n1023, n1027, n1032, n1037, n1042, n1047, n1052, n1057,
    n1062, n1067, n1072, n1077, n1082, n1087, n1092, n1097, n1102, n1107,
    n1112, n1117, n1122, n1127, n1132, n1137, n1142, n1147, n1152, n1157,
    n1162, n1167, n1172, n1176, n1181, n1186, n1191, n1196, n1201, n1206,
    n1211, n1216, n1221, n1226, n1231, n1236, n1241, n1246, n1251, n1256,
    n1261, n1266, n1271, n1276, n1281, n1285, n1290, n1295, n1300, n1305,
    n1310, n1315, n1320, n1325, n1330, n1335, n1340, n1345, n1350, n1355,
    n1360, n1365, n1370, n1374, n1379, n1384, n1389, n1394, n1399, n1403,
    n1408, n1413, n1418, n1423, n1428, n1433, n1438, n1443, n1448, n1453,
    n1458, n1463, n1468, n1473, n1478, n1483, n1488, n1493, n1498, n1502,
    n1506, n1511, n1516, n1521, n1526, n1531, n1536, n1541, n1546, n1551,
    n1556, n1561, n1566, n1571, n1576, n1581, n1585, n1590, n1595, n1600,
    n1605, n1610, n1615, n1620, n1625, n1630, n1635, n1640, n1645, n1650,
    n1655, n1660, n1665, n1669, n1674, n1679, n1684, n1689, n1694, n1699,
    n1704, n1709, n1714, n1719, n1724, n1729, n1734, n1739, n1744, n1749,
    n1754, n1759, n1764, n1768, n1773, n1778, n1783, n1788, n1793, n1798,
    n1803, n1808, n1813, n1818, n1822, n1827, n1832, n1837, n1842, n1847,
    n1851, n1856, n1860, n1865, n1870, n1875, n1880, n1885, n1890, n1895,
    n1900, n1905, n1910, n1915, n1920, n1925, n1930, n1935, n1940, n1945,
    n1950, n1955, n1960, n1965, n1970, n1975, n1980, n1985, n1990, n1995,
    n2000, n2005, n2010, n2014, n2019, n2024, n2029, n2034, n2039, n2044,
    n2049, n2054, n2059, n2064, n2068, n2073, n2078, n2083, n2088, n2093,
    n2098, n2102, n2107, n2111, n2116, n2121, n2125, n2130, n2135, n2140,
    n2145, n2150, n2155, n2160, n2165, n2170, n2175, n2180, n2185, n2190,
    n2195, n2200, n2205, n2210, n2215, n2220, n2225, n2229, n2234, n2238,
    n2243, n2248, n2252, n2257, n2262, n2267, n2271, n2274, n2279, n2284,
    n2289, n2294, n2298, n2303, n2308, n2313, n2318, n2323, n2328, n2333,
    n2338, n2343, n2348, n2353, n2358, n2363, n2368, n2373, n2378, n2383,
    n2388, n2393, n2398, n2403, n2408, n2413, n2418, n2423, n2428, n2433,
    n2438, n2443, n2448, n2453, n2458, n2463, n2467, n2471, n2475, n2478,
    n2482, n2487, n2492, n2497, n2502, n2507, n2512, n2517, n2522, n2527,
    n2532, n2537, n2542, n2547, n2552, n2557, n2562, n2566, n2571, n2576,
    n2581, n2586, n2591, n2596, n2601, n2606, n2610, n2614, n2619, n2624,
    n2629, n2634, n2638, n2643, n2648, n2653, n2658, n2663, n2668, n2673,
    n2678, n2683, n2688, n2693, n2698, n2703, n2708, n2713, n2718, n2722,
    n2727, n2732, n2737, n2742, n2747, n2752, n2757, n2762, n2767, n2771,
    n2775, n2780, n2784, n2789, n2794, n2799, n2804, n2809, n2814, n2819,
    n2824, n2828, n2833, n2837, n2842, n2847, n2852, n2857, n2862, n2867,
    n2872, n2877, n2882, n2887, n2892, n2896, n2901, n2906, n2911, n2916,
    n2921, n2926, n2931, n2936, n2941, n2945, n2950, n2955, n2960, n2965,
    n2968, n2973, n2978, n2982, n2987, n2991, n2996, n3001, n3006, n3011,
    n3016, n3021, n3026, n3031, n3035, n3039, n3043, n3047, n3052, n3055,
    n3060, n3065, n3069, n3074, n3079, n3084, n3089, n3094, n3099, n3104,
    n3109, n3114, n3119, n3124, n3128, n3133, n3138, n3143, n3148, n3153,
    n3158, n3163, n3168, n3173, n3178, n3183, n3188, n3193, n3198, n3202,
    n3207, n3211, n3215, n3220, n3225, n3230, n3235, n3240, n3245, n3249,
    n3253, n3258, n3263, n3268, n3273, n3278, n3282, n3286, n3290, n3295,
    n3300, n3305, n3310, n3315, n3320, n3325, n3329, n3334, n3338, n3342,
    n3347, n3352, n3356, n3361, n3366, n3371, n3376, n3381, n3386, n3391,
    n3396, n3401, n3405, n3409, n3414, n3419, n3424, n3429, n3434, n3439,
    n3444, n3449, n3454, n3459, n3464, n3468, n3473, n3478, n3482, n3487,
    n3492, n3497, n3502, n3506, n3510, n3515, n3520, n3524, n3529, n3534,
    n3539;
  assign g1006 = n2131 & g43 & ~g1000 & g162;
  assign n2131 = n2132 & ~n2383 & ~g1034 & ~n2965 & ~g979 & ~n2054;
  assign n2132 = ~g971 & ~g962 & ~g972 & ~g970 & ~g969 & ~g963 & ~g966;
  assign n2054 = g984 & ~g979 & g43;
  assign n2965 = g973 & g43 & ~g7103 & ~g7298;
  assign g7103 = ~g1 & ~n2132;
  assign g7298 = ~n2132 & g1;
  assign n2383 = g976 & g43 & ~g7298 & ~g7103;
  assign g1015 = n2139 & g1 & ~g1034 & g162;
  assign n2139 = n2132 & g1013 & ~n2383 & ~n2054 & ~g979 & ~n2965;
  assign g4655 = n2141 | n2142;
  assign n2141 = ~g940 & g936;
  assign n2142 = ~g936 & g940;
  assign g4657 = ~g1372 & ~g1371 & ~g1373 & ~g1374 & ~g1375 & ~g1367 & ~g1368 & ~g1369 & ~g1370 & ~g1363 & ~g1364 & ~g1366 & ~g1365;
  assign g4660 = ~g1391 & g1392;
  assign g4661 = ~g1395 & g1394;
  assign g4663 = ~g1398 & g1397;
  assign g4664 = ~g1401 & g1400;
  assign g5164 = g888 & g889 & g887;
  assign g6236 = g1189 | g16;
  assign g6849 = ~g888 & ~g889 & ~g887 & ~g778 & ~n2151;
  assign n2151 = ~n2173 & ~n2170_1 & ~n2167 & ~n2164 & ~n2161 & ~n2158 & ~n2152 & ~n2155_1;
  assign n2152 = ~n2153 & ~n2154;
  assign n2153 = g891 & g831;
  assign n2154 = ~g891 & ~g831;
  assign n2155_1 = ~n2156 & ~n2157;
  assign n2156 = g843 & g911;
  assign n2157 = ~g843 & ~g911;
  assign n2158 = ~n2159 & ~n2160_1;
  assign n2159 = g834 & g896;
  assign n2160_1 = ~g834 & ~g896;
  assign n2161 = ~n2162 & ~n2163;
  assign n2162 = g846 & g916;
  assign n2163 = ~g846 & ~g916;
  assign n2164 = ~n2165_1 & ~n2166;
  assign n2165_1 = g921 & g849;
  assign n2166 = ~g921 & ~g849;
  assign n2167 = ~n2168 & ~n2169;
  assign n2168 = g837 & g901;
  assign n2169 = ~g837 & ~g901;
  assign n2170_1 = ~n2171 & ~n2172;
  assign n2171 = g852 & g883;
  assign n2172 = ~g852 & ~g883;
  assign n2173 = ~n2174 & ~n2175_1;
  assign n2174 = g906 & g840;
  assign n2175_1 = ~g906 & ~g840;
  assign g7048 = g855 | ~g944;
  assign g7063 = ~g1412 | ~g1405;
  assign g7283 = ~g7 | ~n2179;
  assign n2179 = n2181 & g58 & n2180_1;
  assign n2180_1 = g86 & g52 & g80 & g83;
  assign n2181 = g68 & ~g74 & ~g71 & ~g77;
  assign g7284 = ~g6 | ~n2179;
  assign g7285 = ~g5 | ~n2179;
  assign g7286 = ~g4 | ~n2179;
  assign g7287 = ~g2 | ~n2179;
  assign g7288 = ~g3 | ~n2179;
  assign g7289 = ~g48 | ~n2179;
  assign g7290 = ~g8 | ~n2179;
  assign g7291 = ~g48 | ~n2190_1;
  assign n2190_1 = n2191 & g58 & n2180_1;
  assign n2191 = ~g74 & ~g77 & ~g68 & ~g71;
  assign g7292 = ~g3 | ~n2190_1;
  assign g7293 = ~g2 | ~n2190_1;
  assign g7294 = ~g4 | ~n2190_1;
  assign g7474 = g45 | n2196;
  assign n2196 = ~g62 & ~g65;
  assign g7514 = ~n2054 & g1034;
  assign g8234 = ~g1033 | g1029 | ~g43;
  assign g8872 = n2200_1 | ~g1;
  assign n2200_1 = ~n2201 & n2203;
  assign n2201 = g999 & n2202;
  assign n2202 = g998 & ~g1000 & ~g1;
  assign n2203 = ~n2965 & ~n2054 & ~g1030;
  assign g8958 = n2205_1 | ~g1;
  assign n2205_1 = n2203 & ~n2201 & ~n2206;
  assign n2206 = ~g10 & g8234;
  assign g9128 = n2208 | n2209;
  assign n2208 = ~g32 & g31;
  assign n2209 = g32 & g30;
  assign g9280 = n784 | ~g62;
  assign n784 = n2212 | n2282;
  assign n2212 = ~n2213 & n2279_1;
  assign n2213 = ~n2214 & ~n2255;
  assign n2214 = ~n2215_1 & n2244;
  assign n2215_1 = ~n2243_1 & ~n2242 & ~n2241 & ~n2240 & ~n2230 & ~n2227 & ~n2225_1 & ~n2216 & ~n2221;
  assign n2216 = g49 & n2217;
  assign n2217 = n2219 & n1900 & n2180_1;
  assign n1900 = g44 & ~g41 & ~g42 & ~g45 & ~g55;
  assign n2219 = ~g68 & n2220_1;
  assign n2220_1 = g74 & ~g77 & g71;
  assign n2221 = g746 & n2222;
  assign n2222 = n2223 & n1900 & n2180_1;
  assign n2223 = n2224 & ~g71 & g68;
  assign n2224 = ~g74 & g77;
  assign n2225_1 = g694 & n2226;
  assign n2226 = n1900 & n2180_1 & n2191;
  assign n2227 = g710 & n2228;
  assign n2228 = n2229_1 & n1900 & n2180_1;
  assign n2229_1 = g71 & ~g74 & ~g68 & ~g77;
  assign n2230 = ~n2239 & ~n2236 & ~n2235 & ~n2226 & ~n2217 & ~n2233 & ~n2228 & ~n2222 & ~n2231;
  assign n2231 = n2232 & n1900 & n2180_1;
  assign n2232 = n2224 & ~g68 & ~g71;
  assign n2233 = n2234_1 & n1900 & n2180_1;
  assign n2234_1 = g71 & g68 & ~g77 & ~g74;
  assign n2235 = n1900 & n2180_1 & n2181;
  assign n2236 = g74 & g77 & n2237 & n1900 & ~g68 & ~g71;
  assign n2237 = g80 & n2238_1;
  assign n2238_1 = ~g86 & ~g83 & ~g52;
  assign n2239 = g74 & g77 & n1900 & g68 & ~g71 & n2237;
  assign n2240 = g685 & n2233;
  assign n2241 = g648 & n2235;
  assign n2242 = g471 & n2236;
  assign n2243_1 = g527 & n2239;
  assign n2244 = ~n2254 & ~n2253 & ~n2252_1 & ~n2251 & ~n2250 & ~n2249 & ~n2248_1 & ~n2247 & ~n2245 & ~n2246;
  assign n2245 = n2223 & n2237;
  assign n2246 = n2224 & g71 & n2237 & g68;
  assign n2247 = n2224 & g71 & ~g68 & n2237;
  assign n2248_1 = n2232 & n2237;
  assign n2249 = n2220_1 & n2237 & g68;
  assign n2250 = g74 & n2237 & ~g77 & ~g68 & ~g71;
  assign n2251 = n2219 & n2237;
  assign n2252_1 = g74 & g68 & n2237 & ~g71 & ~g77;
  assign n2253 = n2234_1 & n2237;
  assign n2254 = n2229_1 & n2237;
  assign n2255 = ~n2244 & ~n2256;
  assign n2256 = ~n2277 & ~n2263 & ~n2261 & ~n2257_1 & ~n2259;
  assign n2257_1 = g774 & n2258;
  assign n2258 = n1900 & n2252_1;
  assign n2259 = g766 & n2260;
  assign n2260 = n1900 & n2253;
  assign n2261 = g758 & n2262_1;
  assign n2262_1 = n1900 & n2254;
  assign n2263 = ~n2264 & n2275;
  assign n2264 = ~n2274_1 & ~n2273 & ~n2265 & ~n2272;
  assign n2265 = ~n2271_1 & ~n2270 & ~n2269 & ~n2268 & ~n2266 & ~n2267_1;
  assign n2266 = n1900 & n2245;
  assign n2267_1 = n1900 & n2251;
  assign n2268 = n1900 & n2247;
  assign n2269 = n1900 & n2248_1;
  assign n2270 = n1900 & n2246;
  assign n2271_1 = n1900 & n2249;
  assign n2272 = g48 & n2266;
  assign n2273 = g852 & n2270;
  assign n2274_1 = g855 & n2271_1;
  assign n2275 = n1900 & ~n2276 & n2237;
  assign n2276 = ~n2220_1 & ~n2224;
  assign n2277 = ~n2275 & ~n2258 & ~n2262_1 & ~n2278 & ~n2260;
  assign n2278 = n1900 & n2250;
  assign n2279_1 = ~n2280 & ~n2281;
  assign n2280 = ~g80 & n2238_1;
  assign n2281 = n2237 & ~g71 & ~g77 & ~g74;
  assign n2282 = ~n2279_1 & ~n2283;
  assign n2283 = ~n2318_1 & ~n2316 & ~n2314 & ~n2312 & ~n2310 & ~n2308_1 & ~n2306 & ~n2304 & ~n2302 & ~n2300 & ~n2298_1 & ~n2296 & ~n2294_1 & ~n2292 & ~n2290 & ~n2288 & ~n2284_1 & ~n2286;
  assign n2284_1 = g632 & n2285;
  assign n2285 = n2237 & n1900 & n2181;
  assign n2286 = g613 & n2287;
  assign n2287 = g74 & g77 & g71 & n1900 & ~g68 & n2280;
  assign n2288 = g600 & n2289_1;
  assign n2289_1 = n2280 & g74 & g77 & n1900 & ~g68 & ~g71;
  assign n2290 = g621 & n2291;
  assign n2291 = g74 & g77 & g71 & g68 & n1900 & n2280;
  assign n2292 = g608 & n2293;
  assign n2293 = n2280 & g74 & g77 & n1900 & ~g71 & g68;
  assign n2294_1 = g553 & n2295;
  assign n2295 = n2280 & n2224 & g71 & n1900 & g68;
  assign n2296 = g390 & n2297;
  assign n2297 = n2280 & n1900 & n2232;
  assign n2298_1 = g446 & n2299;
  assign n2299 = n2280 & n1900 & n2223;
  assign n2300 = g185 & n2301;
  assign n2301 = n2280 & n1900 & n2181;
  assign n2302 = g168 & n2303_1;
  assign n2303_1 = n2280 & n1900 & n2191;
  assign n2304 = g110 & n2305;
  assign n2305 = n2280 & n1900 & n2229_1;
  assign n2306 = g142 & n2307;
  assign n2307 = n2280 & n1900 & n2234_1;
  assign n2308_1 = g365 & n2309;
  assign n2309 = n2280 & n2220_1 & n1900 & g68;
  assign n2310 = g309 & n2311;
  assign n2311 = n2280 & n1900 & n2219;
  assign n2312 = g228 & n2313_1;
  assign n2313_1 = n2280 & g74 & n1900 & ~g77 & ~g68 & ~g71;
  assign n2314 = g284 & n2315;
  assign n2315 = n2280 & g74 & g68 & n1900 & ~g71 & ~g77;
  assign n2316 = g624 & n2317;
  assign n2317 = n2237 & n1900 & n2191;
  assign n2318_1 = ~n2317 & ~n2285 & ~n2319 & ~n2315 & ~n2313_1 & ~n2311 & ~n2309 & ~n2307 & ~n2305 & ~n2303_1 & ~n2301 & ~n2293 & ~n2289_1 & ~n2291 & ~n2287;
  assign n2319 = n2280 & n1900 & n2224;
  assign g9297 = n1082 | ~g62;
  assign n1082 = n2322 | n2343_1;
  assign n2322 = ~n2323_1 & n2279_1;
  assign n2323_1 = ~n2324 & ~n2334;
  assign n2324 = ~n2325 & n2244;
  assign n2325 = ~n2333_1 & ~n2332 & ~n2331 & ~n2330 & ~n2230 & ~n2329 & ~n2328_1 & ~n2326 & ~n2327;
  assign n2326 = g757 & n2217;
  assign n2327 = g741 & n2222;
  assign n2328_1 = g698 & n2226;
  assign n2329 = g714 & n2228;
  assign n2330 = g681 & n2233;
  assign n2331 = g647 & n2235;
  assign n2332 = g468 & n2236;
  assign n2333_1 = g524 & n2239;
  assign n2334 = ~n2244 & ~n2335;
  assign n2335 = ~n2342 & ~n2341 & ~n2277 & ~n2336;
  assign n2336 = ~n2337 & n2275;
  assign n2337 = ~n2340 & ~n2339 & ~n2265 & ~n2338_1;
  assign n2338_1 = g3 & n2266;
  assign n2339 = g849 & n2270;
  assign n2340 = g859 & n2271_1;
  assign n2341 = g765 & n2260;
  assign n2342 = g773 & n2258;
  assign n2343_1 = ~n2279_1 & ~n2344;
  assign n2344 = ~n2361 & ~n2318_1 & ~n2360 & ~n2359 & ~n2358_1 & ~n2357 & ~n2356 & ~n2355 & ~n2354 & ~n2353_1 & ~n2352 & ~n2351 & ~n2350 & ~n2349 & ~n2348_1 & ~n2347 & ~n2345 & ~n2346;
  assign n2345 = g623 & n2317;
  assign n2346 = g620 & n2291;
  assign n2347 = g607 & n2293;
  assign n2348_1 = g612 & n2287;
  assign n2349 = g599 & n2289_1;
  assign n2350 = g550 & n2295;
  assign n2351 = g387 & n2297;
  assign n2352 = g443 & n2299;
  assign n2353_1 = g182 & n2301;
  assign n2354 = g162 & n2303_1;
  assign n2355 = g105 & n2305;
  assign n2356 = g138 & n2307;
  assign n2357 = g362 & n2309;
  assign n2358_1 = g306 & n2311;
  assign n2359 = g225 & n2313_1;
  assign n2360 = g281 & n2315;
  assign n2361 = g631 & n2285;
  assign g9299 = n2116 | ~g62;
  assign n2116 = n2364 | n2384;
  assign n2364 = ~n2365 & n2279_1;
  assign n2365 = ~n2366 & ~n2375;
  assign n2366 = ~n2367 & n2244;
  assign n2367 = ~n2374 & ~n2373_1 & ~n2372 & ~n2230 & ~n2371 & ~n2370 & ~n2368_1 & ~n2369;
  assign n2368_1 = g677 & n2233;
  assign n2369 = g652 & n2235;
  assign n2370 = g465 & n2236;
  assign n2371 = g513 & n2239;
  assign n2372 = g756 & n2217;
  assign n2373_1 = g702 & n2226;
  assign n2374 = g718 & n2228;
  assign n2375 = ~n2244 & ~n2376;
  assign n2376 = ~n2383_1 & ~n2382 & ~n2277 & ~n2377;
  assign n2377 = ~n2378_1 & n2275;
  assign n2378_1 = ~n2381 & ~n2380 & ~n2265 & ~n2379;
  assign n2379 = g863 & n2271_1;
  assign n2380 = g846 & n2270;
  assign n2381 = g2 & n2266;
  assign n2382 = g764 & n2260;
  assign n2383_1 = g772 & n2258;
  assign n2384 = ~n2279_1 & ~n2385;
  assign n2385 = ~n2402 & ~n2318_1 & ~n2401 & ~n2400 & ~n2399 & ~n2398_1 & ~n2397 & ~n2396 & ~n2395 & ~n2394 & ~n2393_1 & ~n2392 & ~n2391 & ~n2390 & ~n2389 & ~n2388_1 & ~n2386 & ~n2387;
  assign n2386 = g622 & n2317;
  assign n2387 = g619 & n2291;
  assign n2388_1 = g606 & n2293;
  assign n2389 = g611 & n2287;
  assign n2390 = g598 & n2289_1;
  assign n2391 = g547 & n2295;
  assign n2392 = g384 & n2297;
  assign n2393_1 = g432 & n2299;
  assign n2394 = g181 & n2301;
  assign n2395 = g158 & n2303_1;
  assign n2396 = g100 & n2305;
  assign n2397 = g134 & n2307;
  assign n2398_1 = g351 & n2309;
  assign n2399 = g303 & n2311;
  assign n2400 = g222 & n2313_1;
  assign n2401 = g270 & n2315;
  assign n2402 = g630 & n2285;
  assign g9305 = n600 | ~g62;
  assign n600 = n2405 | n2424;
  assign n2405 = ~n2406 & n2279_1;
  assign n2406 = ~n2407 & ~n2416;
  assign n2407 = ~n2408_1 & n2244;
  assign n2408_1 = ~n2415 & ~n2414 & ~n2413_1 & ~n2230 & ~n2412 & ~n2411 & ~n2409 & ~n2410;
  assign n2409 = g673 & n2233;
  assign n2410 = g645 & n2235;
  assign n2411 = g462 & n2236;
  assign n2412 = g510 & n2239;
  assign n2413_1 = g753 & n2217;
  assign n2414 = g734 & n2228;
  assign n2415 = g722 & n2226;
  assign n2416 = ~n2244 & ~n2417;
  assign n2417 = ~n2420 & ~n2419 & ~n2277 & ~n2418_1;
  assign n2418_1 = g763 & n2260;
  assign n2419 = g771 & n2258;
  assign n2420 = ~n2421 & n2275;
  assign n2421 = ~n2422 & ~n2423_1;
  assign n2422 = g843 & n2270;
  assign n2423_1 = g4 & n2266;
  assign n2424 = ~n2279_1 & ~n2425;
  assign n2425 = ~n2441 & ~n2440 & ~n2439 & ~n2438_1 & ~n2437 & ~n2436 & ~n2435 & ~n2434 & ~n2433_1 & ~n2432 & ~n2431 & ~n2430 & ~n2429 & ~n2428_1 & ~n2427 & ~n2318_1 & ~n2426;
  assign n2426 = g629 & n2285;
  assign n2427 = g618 & n2291;
  assign n2428_1 = g605 & n2293;
  assign n2429 = g610 & n2287;
  assign n2430 = g597 & n2289_1;
  assign n2431 = g573 & n2295;
  assign n2432 = g381 & n2297;
  assign n2433_1 = g429 & n2299;
  assign n2434 = g180 & n2301;
  assign n2435 = g154 & n2303_1;
  assign n2436 = g95 & n2305;
  assign n2437 = g130 & n2307;
  assign n2438_1 = g348 & n2309;
  assign n2439 = g300 & n2311;
  assign n2440 = g219 & n2313_1;
  assign n2441 = g267 & n2315;
  assign g9308 = n864 | ~g62;
  assign n864 = n2444 | n2463_1;
  assign n2444 = ~n2445 & n2279_1;
  assign n2445 = ~n2446 & ~n2455;
  assign n2446 = ~n2447 & n2244;
  assign n2447 = ~n2454 & ~n2453_1 & ~n2452 & ~n2230 & ~n2451 & ~n2450 & ~n2448_1 & ~n2449;
  assign n2448_1 = g669 & n2233;
  assign n2449 = g635 & n2235;
  assign n2450 = g459 & n2236;
  assign n2451 = g507 & n2239;
  assign n2452 = g752 & n2217;
  assign n2453_1 = g723 & n2226;
  assign n2454 = g730 & n2228;
  assign n2455 = ~n2244 & ~n2456;
  assign n2456 = ~n2459 & ~n2458_1 & ~n2277 & ~n2457;
  assign n2457 = g762 & n2260;
  assign n2458_1 = g770 & n2258;
  assign n2459 = ~n2460 & n2275;
  assign n2460 = ~n2461 & ~n2462;
  assign n2461 = g840 & n2270;
  assign n2462 = g5 & n2266;
  assign n2463_1 = ~n2279_1 & ~n2464;
  assign n2464 = ~n2480 & ~n2479 & ~n2478_1 & ~n2477 & ~n2476 & ~n2475_1 & ~n2474 & ~n2473 & ~n2472 & ~n2471_1 & ~n2470 & ~n2469 & ~n2468 & ~n2467_1 & ~n2466 & ~n2318_1 & ~n2465;
  assign n2465 = g628 & n2285;
  assign n2466 = g617 & n2291;
  assign n2467_1 = g604 & n2293;
  assign n2468 = g609 & n2287;
  assign n2469 = g596 & n2289_1;
  assign n2470 = g591 & n2295;
  assign n2471_1 = g378 & n2297;
  assign n2472 = g426 & n2299;
  assign n2473 = g179 & n2301;
  assign n2474 = g174 & n2303_1;
  assign n2475_1 = g89 & n2305;
  assign n2476 = g126 & n2307;
  assign n2477 = g345 & n2309;
  assign n2478_1 = g297 & n2311;
  assign n2479 = g216 & n2313_1;
  assign n2480 = g264 & n2315;
  assign g9310 = n1865 | ~g62;
  assign n1865 = n2483 | n2499;
  assign n2483 = ~n2484 & n2279_1;
  assign n2484 = ~n2485 & ~n2491;
  assign n2485 = ~n2486 & n2244;
  assign n2486 = ~n2490 & ~n2230 & ~n2489 & ~n2487_1 & ~n2488;
  assign n2487_1 = g665 & n2233;
  assign n2488 = g504 & n2239;
  assign n2489 = g634 & n2235;
  assign n2490 = g754 & n2217;
  assign n2491 = ~n2244 & ~n2492_1;
  assign n2492_1 = ~n2495 & ~n2494 & ~n2277 & ~n2493;
  assign n2493 = g761 & n2260;
  assign n2494 = g769 & n2258;
  assign n2495 = ~n2496 & n2275;
  assign n2496 = ~n2497_1 & ~n2498;
  assign n2497_1 = g837 & n2270;
  assign n2498 = g6 & n2266;
  assign n2499 = ~n2279_1 & ~n2500;
  assign n2500 = ~n2510 & ~n2509 & ~n2508 & ~n2507_1 & ~n2506 & ~n2505 & ~n2504 & ~n2503 & ~n2502_1 & ~n2318_1 & ~n2501;
  assign n2501 = g616 & n2291;
  assign n2502_1 = g627 & n2285;
  assign n2503 = g261 & n2315;
  assign n2504 = g184 & n2301;
  assign n2505 = g122 & n2307;
  assign n2506 = g150 & n2303_1;
  assign n2507_1 = g603 & n2293;
  assign n2508 = g588 & n2295;
  assign n2509 = g342 & n2309;
  assign n2510 = g423 & n2299;
  assign g9312 = n3220 | ~g62;
  assign n3220 = n2513 | n2529;
  assign n2513 = ~n2514 & n2279_1;
  assign n2514 = ~n2515 & ~n2521;
  assign n2515 = ~n2516 & n2244;
  assign n2516 = ~n2520 & ~n2230 & ~n2519 & ~n2517_1 & ~n2518;
  assign n2517_1 = g661 & n2233;
  assign n2518 = g501 & n2239;
  assign n2519 = g633 & n2235;
  assign n2520 = g755 & n2217;
  assign n2521 = ~n2244 & ~n2522_1;
  assign n2522_1 = ~n2525 & ~n2524 & ~n2277 & ~n2523;
  assign n2523 = g760 & n2260;
  assign n2524 = g768 & n2258;
  assign n2525 = ~n2526 & n2275;
  assign n2526 = ~n2527_1 & ~n2528;
  assign n2527_1 = g834 & n2270;
  assign n2528 = g7 & n2266;
  assign n2529 = ~n2279_1 & ~n2530;
  assign n2530 = ~n2540 & ~n2539 & ~n2538 & ~n2537_1 & ~n2536 & ~n2535 & ~n2534 & ~n2533 & ~n2532_1 & ~n2318_1 & ~n2531;
  assign n2531 = g615 & n2291;
  assign n2532_1 = g626 & n2285;
  assign n2533 = g258 & n2315;
  assign n2534 = g183 & n2301;
  assign n2535 = g118 & n2307;
  assign n2536 = g173 & n2303_1;
  assign n2537_1 = g602 & n2293;
  assign n2538 = g570 & n2295;
  assign n2539 = g339 & n2309;
  assign n2540 = g420 & n2299;
  assign g9314 = n2175 | ~g62;
  assign n2175 = n2543 | n2559;
  assign n2543 = ~n2544 & n2279_1;
  assign n2544 = ~n2545 & ~n2551;
  assign n2545 = ~n2546 & n2244;
  assign n2546 = ~n2550 & ~n2230 & ~n2549 & ~n2547_1 & ~n2548;
  assign n2547_1 = g706 & n2233;
  assign n2548 = g498 & n2239;
  assign n2549 = g690 & n2235;
  assign n2550 = g751 & n2217;
  assign n2551 = ~n2244 & ~n2552_1;
  assign n2552_1 = ~n2555 & ~n2554 & ~n2277 & ~n2553;
  assign n2553 = g759 & n2260;
  assign n2554 = g767 & n2258;
  assign n2555 = ~n2556 & n2275;
  assign n2556 = ~n2557_1 & ~n2558;
  assign n2557_1 = g831 & n2270;
  assign n2558 = g8 & n2266;
  assign n2559 = ~n2279_1 & ~n2560;
  assign n2560 = ~n2569 & ~n2318_1 & ~n2568 & ~n2567 & ~n2566_1 & ~n2565 & ~n2564 & ~n2563 & ~n2561 & ~n2562_1;
  assign n2561 = g614 & n2291;
  assign n2562_1 = g601 & n2293;
  assign n2563 = g417 & n2299;
  assign n2564 = g563 & n2295;
  assign n2565 = g336 & n2309;
  assign n2566_1 = g255 & n2315;
  assign n2567 = g114 & n2307;
  assign n2568 = g146 & n2303_1;
  assign n2569 = g625 & n2285;
  assign g9378 = n2303 | ~g62;
  assign n2303 = n2572 | n2599;
  assign n2572 = ~g44 & n1870;
  assign n1870 = n2574 | n2598;
  assign n2574 = ~n2575 & ~n2595;
  assign n2575 = ~n2576_1 & ~n2594;
  assign n2576_1 = ~n2577 & ~n2585;
  assign n2577 = ~n2578 & ~n2584;
  assign n2578 = ~n2581_1 & ~n2579 & ~n2580;
  assign n2579 = g8 & g7;
  assign n2580 = ~g8 & ~g7;
  assign n2581_1 = ~n2583 & ~n2582 & ~n2579 & ~n2580;
  assign n2582 = g5 & g6;
  assign n2583 = ~g5 & ~g6;
  assign n2584 = ~n2581_1 & ~n2582 & ~n2583;
  assign n2585 = ~n2577 & ~n2586_1;
  assign n2586_1 = ~n2587 & ~n2593;
  assign n2587 = ~n2590 & ~n2588 & ~n2589;
  assign n2588 = g4 & g2;
  assign n2589 = ~g4 & ~g2;
  assign n2590 = ~n2592 & ~n2591_1 & ~n2588 & ~n2589;
  assign n2591_1 = g48 & g3;
  assign n2592 = ~g48 & ~g3;
  assign n2593 = ~n2590 & ~n2591_1 & ~n2592;
  assign n2594 = ~n2586_1 & ~n2585;
  assign n2595 = ~n2575 & ~n2596_1;
  assign n2596_1 = ~n2597 & g47;
  assign n2597 = ~g45 & g44;
  assign n2598 = ~n2596_1 & ~n2595;
  assign n2599 = g44 & ~n2600 & ~n2618;
  assign n2600 = ~n2601_1 & ~n2609;
  assign n2601_1 = ~n2602 & ~n2608;
  assign n2602 = ~n2605 & ~n2603 & ~n2604;
  assign n2603 = n2116 & n600;
  assign n2604 = ~n2116 & ~n600;
  assign n2605 = ~n2607 & ~n2606_1 & ~n2603 & ~n2604;
  assign n2606_1 = n784 & n1082;
  assign n2607 = ~n784 & ~n1082;
  assign n2608 = ~n2605 & ~n2606_1 & ~n2607;
  assign n2609 = ~n2601_1 & ~n2610_1;
  assign n2610_1 = ~n2611 & ~n2617;
  assign n2611 = ~n2614_1 & ~n2612 & ~n2613;
  assign n2612 = n3220 & n2175;
  assign n2613 = ~n3220 & ~n2175;
  assign n2614_1 = ~n2616 & ~n2615 & ~n2612 & ~n2613;
  assign n2615 = n864 & n1865;
  assign n2616 = ~n864 & ~n1865;
  assign n2617 = ~n2614_1 & ~n2615 & ~n2616;
  assign n2618 = ~n2610_1 & ~n2609;
  assign g7763 = ~n2620 & ~n2625;
  assign n2620 = g786 & n2621;
  assign n2621 = g828 & n2622;
  assign n2622 = g825 & n2623;
  assign n2623 = g822 & n2624_1;
  assign n2624_1 = g819 & g815;
  assign n2625 = ~g786 & ~n2621;
  assign n435 = ~g1034 & g154;
  assign n455 = g8 | ~n2141;
  assign n465 = ~n2629_1 & g190;
  assign n2629_1 = ~g207 & ~n2630;
  assign n2630 = ~n2631 & ~n2632;
  assign n2631 = g1206 & g210;
  assign n2632 = ~g1206 & ~g210;
  assign n470 = n2636 | ~n2634_1;
  assign n2634_1 = ~g1553 & ~n2635;
  assign n2635 = g1528 & g1532 & g1537 & g1541 & g1545 & ~g1251 & g1549;
  assign n2636 = n2634_1 & ~n2637 & ~n2639;
  assign n2637 = ~g1541 & ~n2638_1;
  assign n2638_1 = g1528 & g1532 & ~g1251 & g1537;
  assign n2639 = g1528 & g1532 & g1537 & ~g1251 & g1541;
  assign n475 = n2641 | n2642;
  assign n2641 = g1077 & g1084;
  assign n2642 = g1158 & g1176 & g652;
  assign n480 = ~n2644 & g4655;
  assign n2644 = g945 & n2645;
  assign n2645 = g955 & g959;
  assign n485 = g7298 & ~g7103 & g43;
  assign n490 = n2648_1 | n2649;
  assign n2648_1 = g480 & n2236;
  assign n2649 = ~n2236 & g498;
  assign n500 = ~n2651 & ~n2655;
  assign n2651 = ~n2652 & ~n2654;
  assign n2652 = ~n2653_1 & g1092;
  assign n2653_1 = ~g1251 & g1158;
  assign n2654 = ~g1092 & n2653_1;
  assign n2655 = g1073 & g1158;
  assign n510 = ~n2657 & g190;
  assign n2657 = ~g196 & ~n2658_1;
  assign n2658_1 = ~n2659 & ~n2660;
  assign n2659 = g1194 & g195;
  assign n2660 = ~g1194 & ~g195;
  assign n530 = ~n2662 & ~n2663_1;
  assign n2662 = g608 & g1207;
  assign n2663_1 = ~g608 & ~g1207;
  assign n535 = n2677 | n2676 | n2675 | n2674 | n2673_1 | n2672 | n2671 | n2670 | n2669 | n2668_1 | n2667 | n2665 | n2666;
  assign n2665 = g694 & g710;
  assign n2666 = g698 & g714;
  assign n2667 = g723 & g730;
  assign n2668_1 = g702 & g718;
  assign n2669 = g647 & g681;
  assign n2670 = g690 & g706;
  assign n2671 = g648 & g685;
  assign n2672 = g635 & g669;
  assign n2673_1 = g652 & g677;
  assign n2674 = g645 & g673;
  assign n2675 = g722 & g734;
  assign n2676 = g634 & g665;
  assign n2677 = g633 & g661;
  assign n545 = n2679 | n2681;
  assign n2679 = g355 & n2680;
  assign n2680 = ~g368 & g371;
  assign n2681 = ~n2680 & g359;
  assign n550 = ~n2683_1 & ~n2684;
  assign n2683_1 = g620 & g1211;
  assign n2684 = ~g620 & ~g1211;
  assign n555 = ~n2686 & g1247;
  assign n2686 = ~n2687 & ~n2691;
  assign n2687 = ~g1339 & ~n2688_1;
  assign n2688_1 = ~g1339 & ~n2689;
  assign n2689 = g1336 & n2690;
  assign n2690 = g1333 & g1330;
  assign n2691 = ~n2689 & ~n2688_1;
  assign n560 = n2723 | n2720 | n2717 | n2714 | n2711 | n2708_1 | n2705 | n2702 | n2699 | n2693_1 | n2696;
  assign n2693_1 = ~n2694 & ~n2695;
  assign n2694 = g625 & g1351;
  assign n2695 = ~g625 & ~g1351;
  assign n2696 = ~n2697 & ~n2698_1;
  assign n2697 = g624 & g1354;
  assign n2698_1 = ~g624 & ~g1354;
  assign n2699 = ~n2700 & ~n2701;
  assign n2700 = g623 & g1357;
  assign n2701 = ~g623 & ~g1357;
  assign n2702 = ~n2703_1 & ~n2704;
  assign n2703_1 = g622 & g1360;
  assign n2704 = ~g622 & ~g1360;
  assign n2705 = ~n2706 & ~n2707;
  assign n2706 = g632 & g1330;
  assign n2707 = ~g632 & ~g1330;
  assign n2708_1 = ~n2709 & ~n2710;
  assign n2709 = g631 & g1333;
  assign n2710 = ~g631 & ~g1333;
  assign n2711 = ~n2712 & ~n2713_1;
  assign n2712 = g630 & g1336;
  assign n2713_1 = ~g630 & ~g1336;
  assign n2714 = ~n2715 & ~n2716;
  assign n2715 = g629 & g1339;
  assign n2716 = ~g629 & ~g1339;
  assign n2717 = ~n2718_1 & ~n2719;
  assign n2718_1 = g628 & g1342;
  assign n2719 = ~g628 & ~g1342;
  assign n2720 = ~n2721 & ~n2722_1;
  assign n2721 = g627 & g1345;
  assign n2722_1 = ~g627 & ~g1345;
  assign n2723 = ~n2724 & ~n2725;
  assign n2724 = g626 & g1348;
  assign n2725 = ~g626 & ~g1348;
  assign n580 = n1196 | g1173 | g1167 | g1170 | g1166;
  assign n1196 = g1087 & g1098 & g1102 & g1106 & g1110 & g1114 & g1118 & g1122 & g1142 & g1126;
  assign n595 = n2729 & ~n2739 & ~n2741;
  assign n2729 = ~n2730 & ~n2736;
  assign n2730 = n2732_1 & g1519 & g1472 & g1467 & g1462 & g1499 & ~n2733 & ~n2731 & ~g1251;
  assign n2731 = ~g1034 & g150;
  assign n2732_1 = g1481 & g1494 & g1489;
  assign n2733 = ~n2734 & ~n2735;
  assign n2734 = ~g174 & g1514;
  assign n2735 = g1504 & g174 & g1477;
  assign n2736 = n2731 & ~n2737_1 & ~n2738;
  assign n2737_1 = g1513 & g1524;
  assign n2738 = ~g1513 & ~g1524;
  assign n2739 = ~g1477 & ~n2740;
  assign n2740 = n2732_1 & g1499 & g1504 & g1509 & g1514 & g1519 & g1462 & g1467 & ~g1251 & g1472;
  assign n2741 = n2732_1 & g1499 & g1504 & g1509 & g1514 & g1519 & g1462 & g1467 & g1472 & ~g1251 & g1477;
  assign n614 = n2743 | n2745;
  assign n2743 = g456 & n2744;
  assign n2744 = ~g530 & g533;
  assign n2745 = ~n2744 & g465;
  assign n634 = n2747_1 | n2749;
  assign n2747_1 = g233 & n2748;
  assign n2748 = ~g287 & g290;
  assign n2749 = ~n2748 & g243;
  assign n639 = n2729 & ~n2751 & ~n2753;
  assign n2751 = ~g1499 & ~n2752_1;
  assign n2752_1 = ~g1251 & n2732_1;
  assign n2753 = n2732_1 & ~g1251 & g1499;
  assign n649 = ~g1444 | ~n2755;
  assign n2755 = ~g1459 & ~n2756;
  assign n2756 = g1454 & g1450;
  assign n654 = ~n2758 | g1220 | g1217;
  assign n2758 = g1214 & g1211;
  assign n664 = n2760 | n2761;
  assign n2760 = g405 & n2297;
  assign n2761 = ~n2297 & g423;
  assign n674 = ~n2769 & n2763;
  assign n2763 = ~n2764 & g781;
  assign n2764 = g775 & n2765;
  assign n2765 = g812 & n2766;
  assign n2766 = g809 & n2767_1;
  assign n2767_1 = g806 & n2768;
  assign n2768 = g803 & g799;
  assign n2769 = ~n2770 & n2763;
  assign n2770 = ~n2768 & ~n2771_1;
  assign n2771_1 = ~g803 & ~g799;
  assign n714 = n2965 & ~g979 & g43;
  assign n729 = n2774 | n2775_1;
  assign n2774 = g521 & n2236;
  assign n2775_1 = ~n2236 & g527;
  assign n739 = n2777 | n2778;
  assign n2777 = g274 & n2748;
  assign n2778 = ~n2748 & g278;
  assign n744 = ~n2780_1 & ~n2781;
  assign n2780_1 = g1229 & g610;
  assign n2781 = ~g1229 & ~g610;
  assign n749 = n2783 | n2785;
  assign n2783 = ~n2784_1 & g718;
  assign n2784_1 = n2229_1 & g58 & n2180_1;
  assign n2785 = g2 & n2784_1;
  assign n764 = n2788 | g1304 | n2787;
  assign n2787 = ~g1307 & g1288;
  assign n2788 = ~n2789_1 & g1307;
  assign n2789_1 = ~n3300 & ~n2791;
  assign n3300 = g1276 & g1296 & g1284 & g1280 & g1300 & g1288 & g1272 & g1292;
  assign n2791 = ~n2792 & ~n2796;
  assign n2792 = ~g1288 & ~n2793;
  assign n2793 = g1284 & n2794_1;
  assign n2794_1 = g1280 & n2795;
  assign n2795 = g1276 & g1272;
  assign n2796 = n2795 & g1288 & g1280 & g1284;
  assign n769 = ~n2798 & ~n2799_1;
  assign n2798 = g614 & g1225;
  assign n2799_1 = ~g614 & ~g1225;
  assign n789 = n2801 | n2802;
  assign n2801 = g356 & n2311;
  assign n2802 = ~n2311 & g362;
  assign n799 = n2804_1 | n2805;
  assign n2804_1 = g252 & n2313_1;
  assign n2805 = ~n2313_1 & g270;
  assign n809 = n2807 | n2808;
  assign n2807 = ~n2784_1 & g710;
  assign n2808 = g48 & n2784_1;
  assign n814 = n2810 | n2811;
  assign n2810 = ~n2784_1 & g730;
  assign n2811 = g5 & n2784_1;
  assign n824 = ~n2815 & ~n2655 & ~n2813;
  assign n2813 = ~g1037 & ~n2814_1;
  assign n2814_1 = g1130 & g1092 & g1134 & g1138 & n2653_1 & g1149;
  assign n2815 = g1130 & g1092 & g1134 & g1138 & g1149 & n2653_1 & g1037;
  assign n829 = ~n2819_1 & ~g1097 & ~n2817;
  assign n2817 = ~g1102 & ~n2818;
  assign n2818 = g1087 & g1148 & g1098;
  assign n2819_1 = g1087 & g1098 & g1148 & g1102;
  assign n834 = n2821 | n2822;
  assign n2821 = g475 & n2744;
  assign n2822 = ~n2744 & g483;
  assign n839 = ~n2824_1 & n2763;
  assign n2824_1 = g781 & ~g775 & ~n2765;
  assign n849 = ~n2826 & ~n2827;
  assign n2826 = g598 & g1228;
  assign n2827 = ~g598 & ~g1228;
  assign n854 = ~n2829 & n2755;
  assign n2829 = ~n2830 & ~n2833_1;
  assign n2830 = ~g1454 & ~n2831;
  assign n2831 = ~g1454 & ~n2832;
  assign n2832 = g1444 & g1450;
  assign n2833_1 = ~n2832 & ~n2831;
  assign n859 = ~n2838 & ~g1304 & ~n2835;
  assign n2835 = ~g1296 & ~n2836;
  assign n2836 = g1300 & n2837_1 & g1307;
  assign n2837_1 = g1292 & n2793 & g1288;
  assign n2838 = g1307 & g1296 & g1300 & n2837_1;
  assign n869 = ~n2840 & n2634_1;
  assign n2840 = ~n2841 & ~n2842_1;
  assign n2841 = g1532 & g1251;
  assign n2842_1 = ~g1532 & ~g1251;
  assign n879 = n2844 | n2848;
  assign n2844 = ~n2845 & ~n2847_1;
  assign n2845 = ~g741 & ~n2846;
  assign n2846 = n2303 & ~g44 & ~g45 & ~g41 & ~g741 & ~g42;
  assign n2847_1 = n2223 & g58 & n2180_1;
  assign n2848 = g3 & n2847_1;
  assign n884 = ~g1329 & ~n2850;
  assign n2850 = ~g13 & ~n2851;
  assign n2851 = g1325 & g1324 & g1328 & g1327 & g1326 & n2852_1 & g1313;
  assign n2852_1 = g1321 & g1322 & g1323 & n2853 & g1320 & g1319;
  assign n2853 = g1317 & g1318;
  assign n908 = ~g1431 & ~n2855 & ~g1430;
  assign n2855 = g1412 & g1415;
  assign n913 = n2857_1 | n2858;
  assign n2857_1 = g315 & n2680;
  assign n2858 = ~n2680 & g327;
  assign n918 = n2881 | n2878 | n2875 | n2872_1 | n2869 | n2866 | n2860 | n2863;
  assign n2860 = ~n2861 & ~n2862_1;
  assign n2861 = g767 & g1296;
  assign n2862_1 = ~g767 & ~g1296;
  assign n2863 = ~n2864 & ~n2865;
  assign n2864 = g768 & g1300;
  assign n2865 = ~g768 & ~g1300;
  assign n2866 = ~n2867_1 & ~n2868;
  assign n2867_1 = g1292 & g769;
  assign n2868 = ~g1292 & ~g769;
  assign n2869 = ~n2870 & ~n2871;
  assign n2870 = g1288 & g770;
  assign n2871 = ~g1288 & ~g770;
  assign n2872_1 = ~n2873 & ~n2874;
  assign n2873 = g771 & g1284;
  assign n2874 = ~g771 & ~g1284;
  assign n2875 = ~n2876 & ~n2877_1;
  assign n2876 = g772 & g1280;
  assign n2877_1 = ~g772 & ~g1280;
  assign n2878 = ~n2879 & ~n2880;
  assign n2879 = g773 & g1276;
  assign n2880 = ~g773 & ~g1276;
  assign n2881 = ~n2882_1 & ~n2883;
  assign n2882_1 = g774 & g1272;
  assign n2883 = ~g774 & ~g1272;
  assign n923 = ~g1385 & ~g1384 & ~g1386 & ~g1387 & ~g1388 & ~g1380 & ~g1381 & ~g1382 & ~g1383 & ~g1377 & ~g1376 & ~g1379 & ~g1378;
  assign n933 = ~n2886 & ~n2887_1;
  assign n2886 = g1211 & g607;
  assign n2887_1 = ~g1211 & ~g607;
  assign n948 = ~g43 & ~n2889;
  assign n2889 = ~n2890 & ~n2893;
  assign n2890 = ~g985 & ~n2891;
  assign n2891 = g995 & n2892_1;
  assign n2892_1 = ~g985 & ~g990;
  assign n2893 = g985 & n2891;
  assign n978 = ~n2897 & ~n2655 & ~n2895;
  assign n2895 = ~g1138 & ~n2896_1;
  assign n2896_1 = g1130 & g1092 & n2653_1 & g1134;
  assign n2897 = g1130 & g1092 & g1134 & n2653_1 & g1138;
  assign n988 = n2910 | n2899 | n2909;
  assign n2899 = ~g926 & ~n2900;
  assign n2900 = ~n2907 & ~n2901_1 & ~n2906_1;
  assign n2901_1 = ~n2904 & ~n2799 & ~g888 & ~g887 & ~g889;
  assign n2799 = g871 & n2903;
  assign n2903 = g929 & g933;
  assign n2904 = ~g866 & ~n2905;
  assign n2905 = ~g916 & ~g911 & ~g921 & ~g883 & ~g896 & ~g891 & ~g906 & ~g901;
  assign n2906_1 = g889 & ~g887 & ~g888;
  assign n2907 = ~g866 & n2908;
  assign n2908 = g888 & g887 & ~g875 & ~g889;
  assign n2909 = g888 & g889 & ~n2799 & g887;
  assign n2910 = g874 & g889 & ~g888 & g887;
  assign n993 = n2912 | n2914;
  assign n2912 = g377 & n2913;
  assign n2913 = ~g449 & g452;
  assign n2914 = ~n2913 & g390;
  assign n1003 = n2916_1 | n2917;
  assign n2916_1 = g399 & n2297;
  assign n2917 = ~n2297 & g417;
  assign n1008 = n2919 | n2921_1;
  assign n2919 = ~n2920 & g681;
  assign n2920 = n2234_1 & g58 & n2180_1;
  assign n2921_1 = g3 & n2920;
  assign n1013 = n2923 | n2924;
  assign n2923 = g435 & n2913;
  assign n2924 = ~n2913 & g437;
  assign n1018 = n2926_1 | n2927;
  assign n2926_1 = g333 & n2311;
  assign n2927 = ~n2311 & g351;
  assign n1032 = ~n2931_1 & ~n2655 & ~n2929;
  assign n2929 = ~g1049 & ~n2930;
  assign n2930 = g1130 & g1092 & g1134 & g1138 & g1149 & g1037 & g1041 & n2653_1 & g1045;
  assign n2931_1 = g1130 & g1092 & g1134 & g1138 & g1149 & g1037 & g1041 & g1045 & n2653_1 & g1049;
  assign n1037 = ~n2933 & ~g1097 & ~n2818;
  assign n2933 = ~g1098 & ~n2934;
  assign n2934 = g1087 & g1148;
  assign n1047 = n2936_1 | n2937;
  assign n2936_1 = g232 & n2748;
  assign n2937 = ~n2748 & g240;
  assign n1067 = g1228 | g1227 | g1229 | g1230 | g1223 | g1224 | g1226 | g1225;
  assign n1072 = n2940 | n2941_1;
  assign n2940 = g213 & n2748;
  assign n2941_1 = ~n2748 & g222;
  assign n1077 = n2943 | n2944;
  assign n2943 = g402 & n2297;
  assign n2944 = ~n2297 & g420;
  assign n1097 = n2946 | n2947;
  assign n2946 = g376 & n2913;
  assign n2947 = ~n2913 & g387;
  assign n1107 = n2949 | n2950_1;
  assign n2949 = g359 & n2311;
  assign n2950_1 = ~n2311 & g365;
  assign n1112 = n2952 | n2955_1;
  assign n2952 = ~n2954 & ~n2731 & ~n2953;
  assign n2953 = g1486 & n2730;
  assign n2954 = ~g1486 & ~n2730;
  assign n2955_1 = ~g1524 & n2731;
  assign n1117 = n2729 & ~n2957 & ~n2958;
  assign n2957 = ~g1504 & ~n2753;
  assign n2958 = n2732_1 & g1499 & ~g1251 & g1504;
  assign n1127 = ~n2960_1 & ~n2961;
  assign n2960_1 = g619 & g1214;
  assign n2961 = ~g619 & ~g1214;
  assign n1137 = n2620 | n2963;
  assign n2963 = ~n2623 & ~n2964;
  assign n2964 = ~g822 & ~n2624_1;
  assign n1142 = ~n2968_1 & n2966;
  assign n2966 = ~n2967 & g43;
  assign n2967 = ~g1034 & g8234;
  assign n2968_1 = ~g1029 & ~n2969;
  assign n2969 = ~n2970 & g1025;
  assign n2970 = ~g1018 & ~g1021;
  assign n1157 = n2972 | n2974;
  assign n2972 = ~n2973_1 & g174;
  assign n2973_1 = n2280 & g58 & n2191;
  assign n2974 = g5 & n2973_1;
  assign n1162 = n2976 | n2977;
  assign n2976 = ~n2920 & g685;
  assign n2977 = g48 & n2920;
  assign n1167 = ~n2979 & ~g1097 & ~n2934;
  assign n2979 = ~g1087 & ~g1148;
  assign n1181 = n2986 | g1231 | n2981;
  assign n2981 = ~n2982_1 & ~n2985;
  assign n2982_1 = g1207 & n2983;
  assign n2983 = n2984 & n2758 & g1220 & g1217;
  assign n2984 = g1223 & g1225 & g1224;
  assign n2985 = ~g1226 & ~n2982_1;
  assign n2986 = ~g1226 & ~n2985;
  assign n1191 = ~n2988 & ~n2655 & ~n2930;
  assign n2988 = ~g1045 & ~n2989;
  assign n2989 = g1130 & g1092 & g1134 & g1138 & g1149 & g1037 & n2653_1 & g1041;
  assign n1201 = ~n2991_1 & ~n2992;
  assign n2991_1 = g1217 & g605;
  assign n2992 = ~g1217 & ~g605;
  assign n1216 = ~n2645 & ~n2994;
  assign n2994 = ~g959 & ~n2995;
  assign n2995 = ~g959 & g955;
  assign n1221 = ~n2997 & ~n2998;
  assign n2997 = g1225 & g601;
  assign n2998 = ~g1225 & ~g601;
  assign n1226 = n3000 & n2139 & ~g1034 & ~g162;
  assign n3000 = g1 & g43 & g10;
  assign n1241 = n3002 | n3003;
  assign n3002 = g474 & n2744;
  assign n3003 = ~n2744 & g480;
  assign n1256 = n3009 | g1443 | n3005;
  assign n3005 = ~n3008 & n3006_1;
  assign n3006_1 = ~g33 & n3007;
  assign n3007 = g1432 & g1439;
  assign n3008 = g38 & n3006_1;
  assign n3009 = ~n3008 & g38;
  assign n1266 = g1431 | g1412 | g1430;
  assign n1271 = n3015 | g1231 | n3012;
  assign n3012 = ~n3013 & ~n3014;
  assign n3013 = n2983 & g1207 & g1226;
  assign n3014 = ~g1227 & ~n3013;
  assign n3015 = ~g1227 & ~n3014;
  assign n1276 = n3017 | n3018;
  assign n3017 = g234 & n2748;
  assign n3018 = ~n2748 & g246;
  assign n1305 = n3020 | n3021_1;
  assign n3020 = g278 & n2313_1;
  assign n3021_1 = ~n2313_1 & g284;
  assign n1315 = n3023 | n3024;
  assign n3023 = g212 & n2748;
  assign n3024 = ~n2748 & g219;
  assign n1320 = n3026_1 | n3027;
  assign n3026_1 = g408 & n2297;
  assign n3027 = ~n2297 & g426;
  assign n1325 = ~n3029 & ~n3030;
  assign n3029 = g621 & g1207;
  assign n3030 = ~g621 & ~g1207;
  assign n1330 = n3032 | ~n2763;
  assign n3032 = ~n2767_1 & ~n3033;
  assign n3033 = ~g806 & ~n2768;
  assign n1350 = g1034 & ~g8234 & ~g146;
  assign n1365 = ~g1263 | ~n3036;
  assign n3036 = g1228 & g1227 & g1226 & g1230 & ~g1229 & n2984;
  assign n1370 = n3038 | n3039_1;
  assign n3038 = ~n2920 & g669;
  assign n3039_1 = g5 & n2920;
  assign n1384 = n3041 | n3042;
  assign n3041 = g214 & n2748;
  assign n3042 = ~n2748 & g225;
  assign n1389 = n3044 | n3045;
  assign n3044 = g275 & n2313_1;
  assign n3045 = ~n2313_1 & g281;
  assign n1394 = ~n2620 & ~n3047_1;
  assign n3047_1 = ~n2620 & ~n3048;
  assign n3048 = ~n2624_1 & ~n3049;
  assign n3049 = ~g819 & ~g815;
  assign n1399 = g1236 | n435;
  assign n1413 = n3055_1 | g1231 | n3052_1;
  assign n3052_1 = ~n3053 & ~n3054;
  assign n3053 = g1207 & n2758;
  assign n3054 = ~g1217 & ~n3053;
  assign n3055_1 = ~g1217 & ~n3054;
  assign n1423 = ~n3057 & ~n3058;
  assign n3057 = g1229 & g597;
  assign n3058 = ~g1229 & ~g597;
  assign n1428 = n2620 | n3060_1;
  assign n3060_1 = ~n2622 & ~n3061;
  assign n3061 = ~g825 & ~n2623;
  assign n1433 = g1247 & ~n2690 & ~n3063;
  assign n3063 = ~g1333 & ~g1330;
  assign n1453 = n2729 & ~n3065_1 & ~n3066;
  assign n3065_1 = ~g1509 & ~n2958;
  assign n3066 = n2732_1 & g1499 & g1504 & ~g1251 & g1509;
  assign n1463 = ~n3068 & n2966;
  assign n3068 = ~g1029 & ~n3069_1;
  assign n3069_1 = ~g1018 & ~n3070;
  assign n3070 = ~g1025 & ~g1021;
  assign n1468 = n3072 | n3073;
  assign n3072 = g580 & n2297;
  assign n3073 = ~n2297 & g588;
  assign n1473 = n2729 & ~n3075 & ~n3077;
  assign n3075 = ~g1467 & ~n3076;
  assign n3076 = n2732_1 & g1499 & g1504 & g1509 & g1514 & g1519 & ~g1251 & g1462;
  assign n3077 = n2732_1 & g1499 & g1504 & g1509 & g1514 & g1519 & g1462 & ~g1251 & g1467;
  assign n1488 = n3079_1 | n3080;
  assign n3079_1 = g476 & n2744;
  assign n3080 = ~n2744 & g486;
  assign n1493 = n3082 | n3083;
  assign n3082 = g458 & n2744;
  assign n3083 = ~n2744 & g471;
  assign n1498 = ~n3085 & ~n3086;
  assign n3085 = g615 & g1224;
  assign n3086 = ~g615 & ~g1224;
  assign n1506 = n3088 | n3089_1;
  assign n3088 = g495 & n2236;
  assign n3089_1 = ~n2236 & g513;
  assign n1521 = n2966 & ~n3092 & ~g1029 & ~n3091;
  assign n3091 = ~g1018 & n3070;
  assign n3092 = ~n2970 & ~n3093;
  assign n3093 = g1018 & g1021;
  assign n1526 = g1416 & ~g1424 & ~g1421;
  assign n1531 = n3096 | n3097;
  assign n3096 = ~n2141 & g951;
  assign n3097 = g4 & n2141;
  assign n1536 = n3100 & g1214 & n3099_1;
  assign n3099_1 = ~g1207 & g1211;
  assign n3100 = g1217 & g1220;
  assign n1541 = n3102 | n3104_1;
  assign n3102 = g579 & n3103;
  assign n3103 = ~g576 & g595;
  assign n3104_1 = ~n3103 & g580;
  assign n1551 = n3106 & n3100 & g1214;
  assign n3106 = ~g1211 & g1207;
  assign n1561 = n3108 | n3109_1;
  assign n3108 = g394 & n2913;
  assign n3109_1 = ~n2913 & g402;
  assign n1571 = ~n3111 & ~n2655 & ~n2989;
  assign n3111 = ~g1041 & ~n2815;
  assign n1576 = n3113 | n3114_1;
  assign n3113 = g292 & n2680;
  assign n3114_1 = ~n2680 & g297;
  assign n1581 = n3116 | n3117;
  assign n3116 = ~n2141 & g953;
  assign n3117 = g3 & n2141;
  assign n1600 = ~n3119_1 & ~n3120;
  assign n3119_1 = g1224 & g602;
  assign n3120 = ~g1224 & ~g602;
  assign n1610 = ~n3122 & ~g43 & ~n2892_1;
  assign n3122 = g985 & g990;
  assign n1620 = n3124_1 | g1443 | n3006_1;
  assign n3124_1 = ~n3007 & g33;
  assign n1625 = n3126 | n3127;
  assign n3126 = ~n2141 & g950;
  assign n3127 = g5 & n2141;
  assign n1630 = ~g799 & n2763;
  assign n1635 = ~n3130 & n2763;
  assign n3130 = ~n3131 & n2763;
  assign n3131 = ~n2765 & ~n3132;
  assign n3132 = ~g812 & ~n2766;
  assign n1640 = n3134 | n3135;
  assign n3134 = g566 & n3103;
  assign n3135 = ~n3103 & g567;
  assign n1650 = n3137 | n3138_1;
  assign n3137 = g317 & n2680;
  assign n3138_1 = ~n2680 & g333;
  assign n1655 = n3140 | n3141;
  assign n3140 = ~n2973_1 & g168;
  assign n3141 = g48 & n2973_1;
  assign n1674 = g1097 | n3143_1;
  assign n3143_1 = ~n3146 & ~g1097 & ~n3144;
  assign n3144 = ~g1126 & ~n3145;
  assign n3145 = g1087 & g1098 & g1102 & g1106 & g1110 & g1114 & g1118 & g1148 & g1122;
  assign n3146 = g1087 & g1098 & g1102 & g1106 & g1110 & g1114 & g1118 & g1122 & g1148 & g1126;
  assign n1684 = n3148_1 | n3149;
  assign n3148_1 = g103 & g1329;
  assign n3149 = ~g1329 & ~n3150;
  assign n3150 = ~n3151 & ~n3154;
  assign n3151 = ~n3152 & ~n3153_1;
  assign n3152 = g1325 & g1324 & g1313 & n2852_1;
  assign n3153_1 = ~g1326 & ~n3152;
  assign n3154 = ~g1326 & ~n3153_1;
  assign n1694 = n3156 | n3157;
  assign n3156 = g296 & n2680;
  assign n3157 = ~n2680 & g309;
  assign n1714 = n3159 | n3160;
  assign n3159 = g556 & n3103;
  assign n3160 = ~n3103 & g557;
  assign n1719 = ~n3162 & ~n3163_1;
  assign n3162 = g1226 & g613;
  assign n3163_1 = ~g1226 & ~g613;
  assign n1724 = n3169 | g1231 | n3165;
  assign n3165 = ~n3166 & ~n3168_1;
  assign n3166 = n3167 & g1217 & g1214;
  assign n3167 = g1207 & g1211;
  assign n3168_1 = ~g1220 & ~n3166;
  assign n3169 = ~g1220 & ~n3168_1;
  assign n1729 = n3171 | n3172;
  assign n3171 = ~n2973_1 & g158;
  assign n3172 = g2 & n2973_1;
  assign n1739 = n3174 | n3175;
  assign n3174 = ~n2920 & g661;
  assign n3175 = g7 & n2920;
  assign n1754 = n3177 | n3178_1;
  assign n3177 = g98 & g1329;
  assign n3178_1 = ~g1329 & ~n3179;
  assign n3179 = ~n3180 & ~n3183_1;
  assign n3180 = ~n3181 & ~n3182;
  assign n3181 = g1325 & g1324 & n2852_1 & g1313 & g1326;
  assign n3182 = ~g1327 & ~n3181;
  assign n3183_1 = ~g1327 & ~n3182;
  assign n1773 = n3185 | n3186;
  assign n3185 = ~n2973_1 & g150;
  assign n3186 = g6 & n2973_1;
  assign n1783 = n3188_1 | n3190;
  assign n3188_1 = ~n3189 & g859;
  assign n3189 = g58 & n2249;
  assign n3190 = g3 & n3189;
  assign n1793 = n3192 | n3193_1;
  assign n3192 = g516 & n2744;
  assign n3193_1 = ~n2744 & g518;
  assign n1798 = n2729 & ~n2740 & ~n3195;
  assign n3195 = ~g1472 & ~n3077;
  assign n1813 = n3197 | n3198_1;
  assign n3197 = g395 & n2913;
  assign n3198_1 = ~n2913 & g405;
  assign n1818 = ~n2891 & ~n3200;
  assign n3200 = ~g1034 & n3201;
  assign n3201 = ~n3202_1 & ~n2201 & ~n2965;
  assign n3202_1 = g1007 & n3000 & ~g1008 & ~g1016;
  assign n1837 = n3204 | n3205;
  assign n3204 = g557 & n2297;
  assign n3205 = ~n2297 & g563;
  assign n1842 = n3207_1 | n3208;
  assign n3207_1 = g492 & n2236;
  assign n3208 = ~n2236 & g510;
  assign n1875 = n3210 | n3211_1;
  assign n3210 = g141 & g1329;
  assign n3211_1 = ~n3213 & ~g1329 & ~n3212;
  assign n3212 = ~g1317 & ~g1313;
  assign n3213 = g1317 & g1313;
  assign n1880 = n3215_1 | n3216;
  assign n3215_1 = g486 & n2236;
  assign n3216 = ~n2236 & g504;
  assign n1885 = n3218 | n3219;
  assign n3218 = ~n2920 & g665;
  assign n3219 = g6 & n2920;
  assign n1890 = n3221 | n3222;
  assign n3221 = g543 & n3103;
  assign n3222 = ~n3103 & g544;
  assign n1905 = ~n3224 & ~n3226;
  assign n3224 = ~g792 & ~n3225_1;
  assign n3225_1 = ~g792 & g795;
  assign n3226 = g795 & g792;
  assign n1910 = n3228 | n3229;
  assign n3228 = g457 & n2744;
  assign n3229 = ~n2744 & g468;
  assign n1915 = ~g815 & ~n2620;
  assign n1920 = ~g1454 & n3232;
  assign n3232 = ~g1444 & g1450;
  assign n1925 = n3234 | n3235_1;
  assign n3234 = g544 & n2297;
  assign n3235_1 = ~n2297 & g553;
  assign n1935 = n3237 | n3238;
  assign n3237 = g483 & n2236;
  assign n3238 = ~n2236 & g501;
  assign n1940 = ~n3240_1 & g1247;
  assign n3240_1 = ~n3241 & ~n3248;
  assign n3241 = ~g1190 & ~n3242;
  assign n3242 = ~g1190 & ~n3243;
  assign n3243 = g1360 & n3244;
  assign n3244 = g1354 & n3245_1 & g1357;
  assign n3245_1 = n3246 & g1351 & g1345 & g1348;
  assign n3246 = g1342 & n3247;
  assign n3247 = g1336 & n2690 & g1339;
  assign n3248 = ~n3243 & ~n3242;
  assign n1960 = n3250 | n3251;
  assign n3250 = g312 & n2680;
  assign n3251 = ~n2680 & g318;
  assign n1970 = n3253_1 | n3254;
  assign n3253_1 = g324 & n2311;
  assign n3254 = ~n2311 & g342;
  assign n1975 = n3099 | ~g1253;
  assign n3099 = ~n3257 & g1247;
  assign n3257 = ~n3258_1 & n3036;
  assign n3258_1 = ~g1263 & ~g1257;
  assign n1985 = ~n3260 & ~n3261;
  assign n3260 = g1227 & g599;
  assign n3261 = ~g1227 & ~g599;
  assign n1990 = ~n3264 & n3263_1;
  assign n3263_1 = ~g1443 & ~n3007;
  assign n3264 = ~n3265 & ~n3268_1;
  assign n3265 = ~g1432 & ~n3266;
  assign n3266 = ~g1432 & ~n3267;
  assign n3267 = g1439 & g1435;
  assign n3268_1 = ~n3267 & ~n3266;
  assign n1995 = ~n3271 & ~n2655 & ~n3270;
  assign n3270 = ~g1053 & ~n2931_1;
  assign n3271 = g1130 & g1092 & g1134 & g1138 & g1149 & g1037 & g1041 & g1045 & g1049 & n2653_1 & g1053;
  assign n2000 = n3273_1 | n3274;
  assign n3273_1 = g236 & n2748;
  assign n3274 = ~n2748 & g252;
  assign n2005 = n3276 | n3277;
  assign n3276 = g316 & n2680;
  assign n3277 = ~n2680 & g330;
  assign n2010 = n3279 | n3280;
  assign n3279 = g246 & n2313_1;
  assign n3280 = ~n2313_1 & g264;
  assign n2019 = ~n3282_1 & g1247;
  assign n3282_1 = ~n3283 & ~n3286_1;
  assign n3283 = ~g1357 & ~n3284;
  assign n3284 = ~g1357 & ~n3285;
  assign n3285 = g1354 & n3245_1;
  assign n3286_1 = ~n3285 & ~n3284;
  assign n2039 = n3288 | n3289;
  assign n3288 = g243 & n2313_1;
  assign n3289 = ~n2313_1 & g261;
  assign n2049 = n3291 | n3292;
  assign n3291 = g535 & n3103;
  assign n3292 = ~n3103 & g536;
  assign n2059 = n3294 | n3295_1;
  assign n3294 = ~n2764 & g778;
  assign n3295_1 = ~g778 & n2764;
  assign n2068 = ~n3299 & ~g1304 & ~n3297;
  assign n3297 = ~g1292 & ~n3298;
  assign n3298 = g1307 & n2793 & g1288;
  assign n3299 = g1307 & g1292 & g1288 & n2793;
  assign n2078 = n3301 | n3304;
  assign n3301 = ~g1084 & ~n3302;
  assign n3302 = ~n3303 & ~g1084 & ~n2641;
  assign n3303 = g1158 & g1179 & g652;
  assign n3304 = ~n3302 & ~n2641 & ~n3303;
  assign n2083 = n3263_1 & ~n3267 & ~n3306;
  assign n3306 = ~g1439 & ~g1435;
  assign n2093 = ~n3310_1 & ~g1304 & ~n3308;
  assign n3308 = ~g1276 & ~n3309;
  assign n3309 = g1307 & g1272;
  assign n3310_1 = g1307 & n2795;
  assign n2098 = n3312 | n3313;
  assign n3312 = ~g859 & g11;
  assign n3313 = g859 & g12;
  assign n2102 = ~g162 & g43;
  assign n2125 = n3316 | n3317;
  assign n3316 = g587 & n3103;
  assign n3317 = ~n3103 & g560;
  assign n2130 = n3322 | g1231 | n3319;
  assign n3319 = ~n3320_1 & ~n3321;
  assign n3320_1 = g1223 & g1220 & n2758 & g1207 & g1217;
  assign n3321 = ~g1224 & ~n3320_1;
  assign n3322 = ~g1224 & ~n3321;
  assign n2135 = n3324 | n3325_1;
  assign n3324 = g129 & g1329;
  assign n3325_1 = ~g1329 & ~n3326;
  assign n3326 = ~n3327 & ~n3330;
  assign n3327 = ~n3328 & ~n3329_1;
  assign n3328 = g1318 & n3213 & g1319;
  assign n3329_1 = ~g1320 & ~n3328;
  assign n3330 = ~g1320 & ~n3329_1;
  assign n2150 = n3332 | n3333;
  assign n3332 = g318 & n2311;
  assign n3333 = ~n2311 & g336;
  assign n2155 = ~n2903 & ~n3335;
  assign n3335 = ~g933 & ~n3336;
  assign n3336 = ~g933 & g929;
  assign n2165 = n3338_1 | n3339;
  assign n3338_1 = g327 & n2311;
  assign n3339 = ~n2311 & g345;
  assign n2180 = ~n3341 & ~n3344;
  assign n3341 = ~n3342_1 & g888;
  assign n3342_1 = ~n3343 & g887;
  assign n3343 = g889 & n2799;
  assign n3344 = ~g887 & ~n3345;
  assign n3345 = ~n3346 & ~n3348;
  assign n3346 = ~g926 & ~n3347_1;
  assign n3347_1 = g866 & ~n2905 & ~g889;
  assign n3348 = ~g889 & n2799;
  assign n2185 = n3350 | n3351;
  assign n3350 = ~n2620 & g789;
  assign n3351 = ~g789 & n2620;
  assign n2190 = n3353 | n3354;
  assign n3353 = ~n2973_1 & g173;
  assign n3354 = g7 & n2973_1;
  assign n2195 = n3356_1 | n3357;
  assign n3356_1 = g540 & n2297;
  assign n3357 = ~n2297 & g550;
  assign n2200 = n3359 | n3360;
  assign n3359 = g237 & n2313_1;
  assign n3360 = ~n2313_1 & g255;
  assign n2205 = n3362 | n3363;
  assign n3362 = ~n2141 & g948;
  assign n3363 = g7 & n2141;
  assign n2220 = ~g1435 | ~n3263_1;
  assign n2238 = n3366_1 | n3367;
  assign n3366_1 = ~n3189 & g855;
  assign n3367 = g48 & n3189;
  assign n2243 = g1254 & ~n3370 & ~g1231 & ~n3369;
  assign n3369 = ~g1214 & ~n3167;
  assign n3370 = g1214 & n3167;
  assign n2248 = g1097 | n3372;
  assign n3372 = ~n3375 & ~g1097 & ~n3373;
  assign n3373 = ~g1110 & ~n3374;
  assign n3374 = g1087 & g1098 & g1102 & g1148 & g1106;
  assign n3375 = g1087 & g1098 & g1102 & g1106 & g1148 & g1110;
  assign n2267 = ~n3063 | n3401_1 | n3398 | n3395 | n3392 | n3389 | n3386_1 | n3383 | n3377 | n3380;
  assign n3377 = ~n3378 & ~n3379;
  assign n3378 = g761 & g1351;
  assign n3379 = ~g761 & ~g1351;
  assign n3380 = ~n3381_1 & ~n3382;
  assign n3381_1 = g760 & g1354;
  assign n3382 = ~g760 & ~g1354;
  assign n3383 = ~n3384 & ~n3385;
  assign n3384 = g1357 & g759;
  assign n3385 = ~g1357 & ~g759;
  assign n3386_1 = ~n3387 & ~n3388;
  assign n3387 = g758 & g1360;
  assign n3388 = ~g758 & ~g1360;
  assign n3389 = ~n3390 & ~n3391_1;
  assign n3390 = g766 & g1336;
  assign n3391_1 = ~g766 & ~g1336;
  assign n3392 = ~n3393 & ~n3394;
  assign n3393 = g1339 & g765;
  assign n3394 = ~g1339 & ~g765;
  assign n3395 = ~n3396_1 & ~n3397;
  assign n3396_1 = g1342 & g764;
  assign n3397 = ~g1342 & ~g764;
  assign n3398 = ~n3399 & ~n3400;
  assign n3399 = g763 & g1345;
  assign n3400 = ~g763 & ~g1345;
  assign n3401_1 = ~n3402 & ~n3403;
  assign n3402 = g762 & g1348;
  assign n3403 = ~g762 & ~g1348;
  assign n2294 = n2729 & ~n3405_1 & ~n3407;
  assign n3405_1 = ~g1489 & ~n3406;
  assign n3406 = ~g1251 & g1481;
  assign n3407 = g1481 & ~g1251 & g1489;
  assign n2323 = ~g1257 | ~n3036;
  assign n2333 = n3410 | n3411;
  assign n3410 = ~g1416 & g7063;
  assign n3411 = g1409 & g1416;
  assign n2343 = g1254 & ~g1231 & ~n3413;
  assign n3413 = ~n3414_1 & ~n3418;
  assign n3414_1 = ~n3415 & ~n3417;
  assign n3415 = n3416 & g1207 & g1228;
  assign n3416 = g1227 & n2983 & g1226;
  assign n3417 = ~g1229 & ~n3415;
  assign n3418 = ~g1229 & ~n3417;
  assign n2348 = n3420 | n3421;
  assign n3420 = ~n3226 & g782;
  assign n3421 = ~g782 & n3226;
  assign n2353 = n3423 | n3424_1;
  assign n3423 = g231 & n2748;
  assign n3424_1 = ~n2748 & g237;
  assign n2363 = n3426 | n3427;
  assign n3426 = g215 & n2748;
  assign n3427 = ~n2748 & g228;
  assign n2368 = n3429_1 | n3430;
  assign n3429_1 = ~n2920 & g706;
  assign n3430 = g8 & n2920;
  assign n2373 = n3432 | n3435;
  assign n3432 = ~n2847_1 & ~n3433;
  assign n3433 = ~g746 & ~n3434_1;
  assign n3434_1 = g55 & ~g42 & ~g41 & ~g45;
  assign n3435 = g48 & n2847_1;
  assign n2378 = n2729 & ~n3076 & ~n3437;
  assign n3437 = ~g1462 & ~n3438;
  assign n3438 = n2732_1 & g1499 & g1504 & g1509 & g1514 & ~g1251 & g1519;
  assign n2408 = n3440 | n3441;
  assign n3440 = ~n2622 & g828;
  assign n3441 = ~g828 & n2622;
  assign n2418 = n3443 | n3444_1;
  assign n3443 = g478 & n2744;
  assign n3444_1 = ~n2744 & g492;
  assign n2428 = n2141 | n3446;
  assign n3446 = ~g943 & g4655;
  assign n2448 = n3448 | n3449_1;
  assign n3448 = g354 & n2680;
  assign n3449_1 = ~n2680 & g356;
  assign n2453 = n3451 | n3452;
  assign n3451 = ~n2141 & g952;
  assign n3452 = g2 & n2141;
  assign n2458 = g1186 | g1182 | g1179 | g1073 | g1160 | g1163;
  assign n2463 = ~n3455 & ~n3456;
  assign n3455 = g612 & g1227;
  assign n3456 = ~g612 & ~g1227;
  assign n2471 = ~g1428 & ~n3458 & ~g1429;
  assign n3458 = g1405 & g1408;
  assign n2482 = n3463 | g1231 | n3460;
  assign n3460 = ~n3461 & ~n3462;
  assign n3461 = g1223 & g1217 & g1224 & n2758 & g1207 & g1220;
  assign n3462 = ~g1225 & ~n3461;
  assign n3463 = ~g1225 & ~n3462;
  assign n2487 = n3465 | n3466;
  assign n3465 = g1130 & g1092 & g1134 & g1138 & g1149 & g1037 & g1041 & g1045 & g1049 & g1053 & g1057 & g1061 & g1065 & g1069 & g1158 & ~g1073 & ~g1251;
  assign n3466 = ~g1158 & g1073;
  assign n2492 = n3468_1 | n3469;
  assign n3468_1 = g113 & g1329;
  assign n3469 = ~g1329 & ~n3470;
  assign n3470 = ~n3471 & ~n3474;
  assign n3471 = ~n3472 & ~n3473_1;
  assign n3472 = g1313 & n2852_1;
  assign n3473_1 = ~g1324 & ~n3472;
  assign n3474 = ~g1324 & ~n3473_1;
  assign n2497 = ~n3478_1 & ~n2655 & ~n3476;
  assign n3476 = ~g1069 & ~n3477;
  assign n3477 = g1130 & g1092 & g1134 & g1138 & g1149 & g1037 & g1041 & g1045 & g1049 & g1053 & g1057 & g1061 & n2653_1 & g1065;
  assign n3478_1 = g1130 & g1092 & g1134 & g1138 & g1149 & g1037 & g1041 & g1045 & g1049 & g1053 & g1057 & g1061 & g1065 & n2653_1 & g1069;
  assign n2502 = n3480 | n3481;
  assign n3480 = g437 & n2297;
  assign n3481 = ~n2297 & g443;
  assign n2507 = ~n3483 & ~n3484;
  assign n3483 = g611 & g1228;
  assign n3484 = ~g611 & ~g1228;
  assign n2552 = n2909 | n2908 | n3486 | n3487_1;
  assign n3486 = g887 & ~g888 & ~g878 & ~g889;
  assign n3487_1 = g866 & n2906_1;
  assign n2557 = n3489 | n3490;
  assign n3489 = g560 & n2297;
  assign n3490 = ~n2297 & g573;
  assign n2562 = n3492_1 | n3493;
  assign n3492_1 = g393 & n2913;
  assign n3493 = ~n2913 & g399;
  assign n2571 = n3495 | n3496;
  assign n3495 = g489 & n2236;
  assign n3496 = ~n2236 & g507;
  assign n2576 = n3498 | n3499;
  assign n3498 = g536 & n2297;
  assign n3499 = ~n2297 & g547;
  assign n2596 = g1231 | ~g1207;
  assign n2601 = n3502_1 | n3503;
  assign n3502_1 = g235 & n2748;
  assign n3503 = ~n2748 & g249;
  assign n2606 = g58 | g65;
  assign n2614 = ~n2142 & g942;
  assign n2629 = ~n2644 & ~n3507;
  assign n3507 = ~g945 & ~n3508;
  assign n3508 = ~g945 & n2645;
  assign n2634 = g1097 | n3510_1;
  assign n3510_1 = ~n3512 & ~g1097 & ~n3511;
  assign n3511 = ~g1114 & ~n3375;
  assign n3512 = g1087 & g1098 & g1102 & g1106 & g1110 & g1148 & g1114;
  assign n2643 = n3514 | n3515_1;
  assign n3514 = g411 & n2297;
  assign n3515_1 = ~n2297 & g429;
  assign n2648 = n3517 | ~n2763;
  assign n3517 = ~n2766 & ~n3518;
  assign n3518 = ~g809 & ~n2767_1;
  assign n2658 = g1428 | g1405 | g1429;
  assign n2663 = g1247 & ~n2689 & ~n3521;
  assign n3521 = ~g1336 & ~n2690;
  assign n2678 = ~n3523 & ~n2655 & ~n3477;
  assign n3523 = ~g1065 & ~n3524_1;
  assign n3524_1 = g1130 & g1092 & g1134 & g1138 & g1149 & g1037 & g1041 & g1045 & g1049 & g1053 & g1057 & n2653_1 & g1061;
  assign n2683 = g1097 | n3526;
  assign n3526 = ~n3145 & ~n3527;
  assign n3527 = ~g1122 & ~n3528;
  assign n3528 = g1087 & g1098 & g1102 & g1106 & g1110 & g1114 & g1148 & g1118;
  assign n2688 = n3533 | g1231 | n3530;
  assign n3530 = ~n3531 & ~n3532;
  assign n3531 = g1207 & n3416;
  assign n3532 = ~g1228 & ~n3531;
  assign n3533 = ~g1228 & ~n3532;
  assign n2693 = n3535 | n3536;
  assign n3535 = g479 & n2744;
  assign n3536 = ~n2744 & g495;
  assign n2698 = n3538 | n3539_1;
  assign n3538 = g121 & g1329;
  assign n3539_1 = ~g1329 & ~n3540;
  assign n3540 = ~n3541 & ~n3544;
  assign n3541 = ~n3542 & ~n3543;
  assign n3542 = g1321 & g1320 & n2853 & g1313 & g1319;
  assign n3543 = ~g1322 & ~n3542;
  assign n3544 = ~g1322 & ~n3543;
  assign n2703 = g1231 | n3546;
  assign n3546 = ~n3547 & g1254;
  assign n3547 = ~n3548 & ~n3551;
  assign n3548 = ~n3549 & ~n3550;
  assign n3549 = g1228 & g1229 & n3013 & g1227;
  assign n3550 = ~g1230 & ~n3549;
  assign n3551 = ~g1230 & ~n3550;
  assign n2708 = ~n2383 & ~n3553;
  assign n3553 = g8234 & ~n3554 & n3201;
  assign n3554 = g1018 & n3070;
  assign n2713 = n3556 | n3557;
  assign n3556 = g249 & n2313_1;
  assign n3557 = ~n2313_1 & g267;
  assign n2737 = g1214 & n3100 & ~g1207 & ~g1211;
  assign n2742 = n3560 | n3561;
  assign n3560 = ~n2784_1 & g714;
  assign n3561 = g3 & n2784_1;
  assign n2747 = n3563 | n3564;
  assign n3563 = ~n2784_1 & g734;
  assign n3564 = g4 & n2784_1;
  assign n2752 = ~n3567 & ~g1097 & ~n3566;
  assign n3566 = ~g1142 & ~n3146;
  assign n3567 = g1148 & n1196;
  assign n2757 = g1247 & ~n3246 & ~n3569;
  assign n3569 = ~g1342 & ~n3247;
  assign n2767 = n3571 | n3572;
  assign n3571 = ~g1176 & g1081;
  assign n3572 = ~g1081 & g1080;
  assign n2771 = n2729 & ~n3406 & ~n3574;
  assign n3574 = ~g1481 & g1251;
  assign n2789 = g1247 & ~n3285 & ~n3576;
  assign n3576 = ~g1354 & ~n3245_1;
  assign n2794 = n3578 | n3579;
  assign n3578 = g477 & n2744;
  assign n3579 = ~n2744 & g489;
  assign n2809 = n3581 | n3582;
  assign n3581 = g584 & n2297;
  assign n3582 = ~n2297 & g591;
  assign n2819 = ~g1269 & ~g1268;
  assign n2842 = n3585 | n3586;
  assign n3585 = ~n2141 & g949;
  assign n3586 = g6 & n2141;
  assign n2852 = n3588 | n3589;
  assign n3588 = g396 & n2913;
  assign n3589 = ~n2913 & g408;
  assign n2857 = ~n2799 & ~n3591;
  assign n3591 = ~g871 & ~n3592;
  assign n3592 = ~g871 & n2903;
  assign n2867 = n3594 | n3595;
  assign n3594 = ~n2973_1 & g146;
  assign n3595 = g8 & n2973_1;
  assign n2872 = ~n3597 & g190;
  assign n3597 = ~g202 & ~n3598;
  assign n3598 = ~n3599 & ~n3600;
  assign n3599 = g1202 & g205;
  assign n3600 = ~g1202 & ~g205;
  assign n2877 = n3602 | n3603;
  assign n3602 = g436 & n2913;
  assign n3603 = ~n2913 & g440;
  assign n2892 = ~n3605 & ~n2655 & ~n2814_1;
  assign n3605 = ~g1149 & ~n2897;
  assign n2916 = n3607 | n3608;
  assign n3607 = g567 & n2297;
  assign n3608 = ~n2297 & g570;
  assign n2921 = n3610 | n3611;
  assign n3610 = g273 & n2748;
  assign n3611 = ~n2748 & g275;
  assign n2926 = n3613 | n3614;
  assign n3613 = g294 & n2680;
  assign n3614 = ~n2680 & g303;
  assign n2950 = n3616 | n3617;
  assign n3616 = g133 & g1329;
  assign n3617 = ~g1329 & ~n3618;
  assign n3618 = ~n3619 & ~n3622;
  assign n3619 = ~n3620 & ~n3621;
  assign n3620 = g1313 & n2853;
  assign n3621 = ~g1319 & ~n3620;
  assign n3622 = ~g1319 & ~n3621;
  assign n2955 = n3624 | n3626;
  assign n3624 = ~n3189 & ~n3625;
  assign n3625 = ~g863 & ~g866;
  assign n3626 = g2 & n3189;
  assign n2960 = n3106 | g1231 | n3099_1;
  assign n2973 = ~n3629 & ~n3630;
  assign n3629 = g1217 & g618;
  assign n3630 = ~g1217 & ~g618;
  assign n2978 = g887 & g878 & ~g889 & g888;
  assign n2987 = ~n3633 & ~n3634;
  assign n3633 = g600 & g1226;
  assign n3634 = ~g600 & ~g1226;
  assign n2996 = n3636 | n3637;
  assign n3636 = g108 & g1329;
  assign n3637 = ~g1329 & ~n3638;
  assign n3638 = ~n3639 & ~n3642;
  assign n3639 = ~n3640 & ~n3641;
  assign n3640 = n2852_1 & g1313 & g1324;
  assign n3641 = ~g1325 & ~n3640;
  assign n3642 = ~g1325 & ~n3641;
  assign n3001 = ~n3645 & ~g1304 & ~n3644;
  assign n3644 = ~g1280 & ~n3310_1;
  assign n3645 = g1307 & n2794_1;
  assign n3006 = g1097 | n3647;
  assign n3647 = ~n3648 & ~g1097 & ~n3374;
  assign n3648 = ~g1106 & ~n2819_1;
  assign n3011 = ~n3650 & ~n2655 & ~n3524_1;
  assign n3650 = ~g1061 & ~n3651;
  assign n3651 = g1130 & g1092 & g1134 & g1138 & g1149 & g1037 & g1041 & g1045 & g1049 & g1053 & n2653_1 & g1057;
  assign n3016 = ~n3653 & ~n3654;
  assign n3653 = g1220 & g617;
  assign n3654 = ~g1220 & ~g617;
  assign n3026 = g1444 & ~g1450 & g1454;
  assign n3031 = n3657 | n3658;
  assign n3657 = g373 & n2913;
  assign n3658 = ~n2913 & g378;
  assign n3039 = n2729 & ~n3660 & ~n3661;
  assign n3660 = ~g1514 & ~n3066;
  assign n3661 = n2732_1 & g1499 & g1504 & g1509 & ~g1251 & g1514;
  assign n3047 = g1247 & ~n3663 & ~n3664;
  assign n3663 = ~g1345 & ~n3246;
  assign n3664 = g1345 & n3246;
  assign n3074 = n3669 | g1231 | n3666;
  assign n3666 = ~n3667 & ~n3668;
  assign n3667 = n2758 & g1217 & g1207 & g1220;
  assign n3668 = ~g1223 & ~n3667;
  assign n3669 = ~g1223 & ~n3668;
  assign n3079 = n3671 | n3672;
  assign n3671 = g440 & n2297;
  assign n3672 = ~n2297 & g446;
  assign n3084 = g1424 | n3674;
  assign n3674 = ~g1421 & ~g1416;
  assign n3104 = n3676 | n3677;
  assign n3676 = g211 & n2748;
  assign n3677 = ~n2748 & g216;
  assign n3119 = n3679 | n3680;
  assign n3679 = g539 & n3103;
  assign n3680 = ~n3103 & g540;
  assign n3128 = n2634_1 & ~n2638_1 & ~n3682;
  assign n3682 = ~g1537 & ~n3683;
  assign n3683 = g1528 & ~g1251 & g1532;
  assign n3133 = n3685 | n3686;
  assign n3685 = ~n2635 & g727;
  assign n3686 = ~g727 & n2635;
  assign n3138 = n2131 & n2202;
  assign n3148 = ~n3689 & ~g1304 & ~n3309;
  assign n3689 = ~g1307 & ~g1272;
  assign n3158 = n3691 | n3692;
  assign n3691 = g93 & g1329;
  assign n3692 = ~g1329 & ~n3693;
  assign n3693 = ~n3694 & ~n3697;
  assign n3694 = ~n3695 & ~n3696;
  assign n3695 = g1327 & g1326 & n3640 & g1325;
  assign n3696 = ~g1328 & ~n3695;
  assign n3697 = ~g1328 & ~n3696;
  assign n3163 = ~n3701 & ~n2655 & ~n3699;
  assign n3699 = ~g1130 & ~n3700;
  assign n3700 = g1092 & n2653_1;
  assign n3701 = g1130 & n2653_1 & g1092;
  assign n3168 = ~g1330 & g1247;
  assign n3188 = n3704 | n3705;
  assign n3704 = g518 & n2236;
  assign n3705 = ~n2236 & g524;
  assign n3193 = ~n3707 & ~n3708;
  assign n3707 = g596 & g1230;
  assign n3708 = ~g596 & ~g1230;
  assign n3198 = n3710 | n3711;
  assign n3710 = g330 & n2311;
  assign n3711 = ~n2311 & g348;
  assign n3207 = g1247 & ~n3713 & ~n3715;
  assign n3713 = ~g1348 & ~n3714;
  assign n3714 = g1345 & n3247 & g1342;
  assign n3715 = g1348 & g1342 & g1345 & n3247;
  assign n3215 = ~g1266 | ~n3036;
  assign n3225 = n3718 | n3719;
  assign n3718 = g240 & n2313_1;
  assign n3719 = ~n2313_1 & g258;
  assign n3230 = n3721 | n3722;
  assign n3721 = g517 & n2744;
  assign n3722 = ~n2744 & g521;
  assign n3235 = n3724 | n3725;
  assign n3724 = g293 & n2680;
  assign n3725 = ~n2680 & g300;
  assign n3245 = g1097 | n3727;
  assign n3727 = ~n3728 & ~g1097 & ~n3528;
  assign n3728 = ~g1118 & ~n3512;
  assign n3253 = n3730 | n3731;
  assign n3730 = g137 & g1329;
  assign n3731 = ~n3733 & ~g1329 & ~n3732;
  assign n3732 = ~g1318 & ~n3213;
  assign n3733 = g1318 & n3213;
  assign n3258 = ~n3735 & ~n3736;
  assign n3735 = g1223 & g603;
  assign n3736 = ~g1223 & ~g603;
  assign n3263 = n3738 | n3739;
  assign n3738 = ~n2920 & g677;
  assign n3739 = g2 & n2920;
  assign n3273 = ~n3741 & ~n2655 & ~n3651;
  assign n3741 = ~g1057 & ~n3271;
  assign n3278 = g7103 & ~g7298 & g43;
  assign n3290 = n2634_1 & ~n2635 & ~n3744;
  assign n3744 = ~g1549 & ~n3745;
  assign n3745 = g1528 & g1532 & g1537 & g1541 & ~g1251 & g1545;
  assign n3295 = n3747 | n3748;
  assign n3747 = g1329 & g125;
  assign n3748 = ~g1329 & ~n3749;
  assign n3749 = ~n3750 & ~n3753;
  assign n3750 = ~n3751 & ~n3752;
  assign n3751 = n2853 & g1319 & g1313 & g1320;
  assign n3752 = ~g1321 & ~n3751;
  assign n3753 = ~g1321 & ~n3752;
  assign n3305 = n2729 & ~n3438 & ~n3755;
  assign n3755 = ~g1519 & ~n3661;
  assign n3310 = n3757 | n3758;
  assign n3757 = g583 & n3103;
  assign n3758 = ~n3103 & g584;
  assign n3320 = n3760 | n3761;
  assign n3760 = g314 & n2680;
  assign n3761 = ~n2680 & g324;
  assign n3325 = n3763 | n3764;
  assign n3763 = g414 & n2297;
  assign n3764 = ~n2297 & g432;
  assign n3334 = n3766 | n3767;
  assign n3766 = g313 & n2680;
  assign n3767 = ~n2680 & g321;
  assign n3342 = n3769 | n3770;
  assign n3769 = g398 & n2913;
  assign n3770 = ~n2913 & g414;
  assign n3347 = ~n3772 & ~n3773;
  assign n3772 = g1220 & g604;
  assign n3773 = ~g1220 & ~g604;
  assign n3356 = ~g1304 & ~n3775;
  assign n3775 = ~n3776 & ~n3777;
  assign n3776 = ~g1307 & g1284;
  assign n3777 = g1307 & ~n3778 & ~n3779;
  assign n3778 = ~g1284 & ~n2794_1;
  assign n3779 = g1284 & g1272 & g1276 & g1280;
  assign n3361 = n3781 | ~n2634_1;
  assign n3781 = n2634_1 & ~n3745 & ~n3782;
  assign n3782 = ~g1545 & ~n2639;
  assign n3366 = ~n3784 & ~n3785;
  assign n3784 = g616 & g1223;
  assign n3785 = ~g616 & ~g1223;
  assign n3371 = n3787 | n3788;
  assign n3787 = ~n2920 & g673;
  assign n3788 = g4 & n2920;
  assign n3381 = n3790 | n3791;
  assign n3790 = g295 & n2680;
  assign n3791 = ~n2680 & g306;
  assign n3386 = n3793 | n3794;
  assign n3793 = ~n2141 & g954;
  assign n3794 = g48 & n2141;
  assign n3391 = n3796 | n3797;
  assign n3796 = ~n2973_1 & g162;
  assign n3797 = g3 & n2973_1;
  assign n3396 = n3799 | n3800;
  assign n3799 = g397 & n2913;
  assign n3800 = ~n2913 & g411;
  assign n3401 = ~g878 & g874;
  assign n3409 = ~n3805 & ~g1304 & ~n3803;
  assign n3803 = ~g1300 & ~n3804;
  assign n3804 = g1307 & n2837_1;
  assign n3805 = n2837_1 & g1307 & g1300;
  assign n3414 = n3807 | n3808;
  assign n3807 = g375 & n2913;
  assign n3808 = ~n2913 & g384;
  assign n3419 = n3810 | n3811;
  assign n3810 = g321 & n2311;
  assign n3811 = ~n2311 & g339;
  assign n3424 = n3813 | n3814;
  assign n3813 = g454 & n2744;
  assign n3814 = ~n2744 & g459;
  assign n3429 = n3816 | n3817;
  assign n3816 = g117 & g1329;
  assign n3817 = ~g1329 & ~n3818;
  assign n3818 = ~n3819 & ~n3822;
  assign n3819 = ~n3820 & ~n3821;
  assign n3820 = g1321 & g1319 & g1322 & n2853 & g1313 & g1320;
  assign n3821 = ~g1323 & ~n3820;
  assign n3822 = ~g1323 & ~n3821;
  assign n3434 = n3824 | n3825;
  assign n3824 = g374 & n2913;
  assign n3825 = ~n2913 & g381;
  assign n3439 = n2634_1 & ~n3683 & ~n3827;
  assign n3827 = ~g1528 & ~n3828;
  assign n3828 = ~g1251 & g1532;
  assign n3444 = ~n3830 & g1247;
  assign n3830 = ~n3831 & ~n3834;
  assign n3831 = ~g1351 & ~n3832;
  assign n3832 = ~g1351 & ~n3833;
  assign n3833 = g1348 & n3714;
  assign n3834 = ~n3833 & ~n3832;
  assign n3454 = ~n3836 & ~n3837;
  assign n3836 = g606 & g1214;
  assign n3837 = ~g606 & ~g1214;
  assign n3459 = ~g172 & ~n3839;
  assign n3839 = ~n3840 & ~n3841;
  assign n3840 = ~n2973_1 & g154;
  assign n3841 = g4 & n2973_1;
  assign n3473 = ~n3843 & ~n2655 & ~n2896_1;
  assign n3843 = ~g1134 & ~n3701;
  assign n3478 = ~n3846 & ~g43 & ~n3845;
  assign n3845 = ~g995 & ~n3122;
  assign n3846 = g995 & n3122;
  assign n3487 = n3848 | n3849;
  assign n3848 = g145 & g1329;
  assign n3849 = ~g1329 & ~g1313;
  assign n3497 = n2729 & ~n2752_1 & ~n3851;
  assign n3851 = ~g1494 & ~n3407;
  assign n3502 = n3853 | n3854;
  assign n3853 = g455 & n2744;
  assign n3854 = ~n2744 & g462;
  assign n3510 = g1247 & ~n3856 & ~n3857;
  assign n3856 = ~g1360 & ~n3244;
  assign n3857 = g1360 & g1354 & g1357 & n3245_1;
  assign n3515 = ~n3859 & n2755;
  assign n3859 = ~n3232 & ~n3860;
  assign n3860 = ~g1450 & g1444;
  assign n3520 = ~n3862 & g190;
  assign n3862 = ~g187 & ~n3863;
  assign n3863 = ~n3864 & ~n3865;
  assign n3864 = g1198 & g186;
  assign n3865 = ~g1198 & ~g186;
  assign n3529 = ~n3867 & ~n3868;
  assign n3867 = g609 & g1230;
  assign n3868 = ~g609 & ~g1230;
  assign g8661 = 1'b0;
  assign n1087 = 1'b0;
  assign g6223 = ~g1486;
  assign g6675 = ~g1432;
  assign g6850 = ~g43;
  assign g6895 = ~g689;
  assign g3856 = ~g929;
  assign g3857 = ~g955;
  assign g3854 = ~g795;
  assign n565 = ~g1260;
  assign n903 = ~g1158;
  assign n1360 = ~g1252;
  assign n2064 = ~g158;
  assign n2308 = ~g1034;
  assign g206 = g1460;
  assign g291 = g1460;
  assign g372 = g1460;
  assign g453 = g1460;
  assign g534 = g1460;
  assign g594 = g1460;
  assign g785 = g888;
  assign g1017 = g1029;
  assign g1246 = g1245;
  assign g1724 = g1409;
  assign g1783 = g891;
  assign g1798 = g921;
  assign g1804 = g916;
  assign g1810 = g911;
  assign g1817 = g906;
  assign g1824 = g901;
  assign g1829 = g896;
  assign g1870 = g963;
  assign g1871 = g966;
  assign g1894 = g1240;
  assign g1911 = g1524;
  assign g1944 = g1081;
  assign g2662 = g1254;
  assign g2844 = g576;
  assign g2888 = g1084;
  assign g3077 = g1029;
  assign g3096 = g287;
  assign g3130 = g368;
  assign g3159 = g449;
  assign g3191 = g530;
  assign g3829 = g1461;
  assign g3859 = g1461;
  assign g3860 = g1461;
  assign g4267 = g1073;
  assign g4316 = g878;
  assign g4370 = g1160;
  assign g4371 = g1163;
  assign g4372 = g1182;
  assign g4373 = g1186;
  assign g5143 = g1554;
  assign g5571 = g1236;
  assign g5669 = g13;
  assign g5678 = g16;
  assign g5682 = g20;
  assign g5684 = g33;
  assign g5687 = g38;
  assign g5729 = g49;
  assign g6207 = g173;
  assign g6212 = g1389;
  assign g6269 = g1000;
  assign g6425 = g1034;
  assign g6648 = g1251;
  assign g6653 = g1250;
  assign g6909 = g1008;
  assign g7295 = g7294;
  assign g7423 = g1167;
  assign g7424 = g1170;
  assign g7425 = g1173;
  assign g7504 = g13;
  assign g7505 = g16;
  assign g7506 = g20;
  assign g7507 = g33;
  assign g7508 = g38;
  assign g7729 = g173;
  assign g7730 = g1389;
  assign g7731 = g6236;
  assign g7732 = ~g1486;
  assign g8216 = g1251;
  assign g8217 = g1250;
  assign g8218 = g1034;
  assign g8219 = ~g1432;
  assign g8663 = g7063;
  assign g9132 = g8234;
  assign g9204 = g9128;
  assign g6294 = g24;
  assign g6376 = g25;
  assign g6300 = g29;
  assign g6292 = g22;
  assign g6298 = g28;
  assign g6291 = g10;
  assign g6293 = g23;
  assign g6304 = g37;
  assign g6296 = g26;
  assign g6289 = g1;
  assign g6297 = g27;
  assign g6306 = g42;
  assign g6290 = g11;
  assign g6303 = g32;
  assign g6305 = g41;
  assign g6302 = g31;
  assign g6308 = g45;
  assign g6288 = g9;
  assign g6307 = g44;
  assign g6299 = g21;
  assign g6301 = g30;
  assign g6295 = g25;
  assign n430 = g1217;
  assign n440 = g1225;
  assign n445 = g1211;
  assign n450 = g449;
  assign n460 = g4;
  assign n495 = g1223;
  assign n505 = g1230;
  assign n515 = g1280;
  assign n520 = g1230;
  assign n525 = g2;
  assign n540 = g10;
  assign n570 = g8;
  assign n575 = g1225;
  assign n585 = g1236;
  assign n590 = g1228;
  assign n605 = g48;
  assign n610 = g1204;
  assign n619 = g48;
  assign n624 = g916;
  assign n629 = g1312;
  assign n644 = g5;
  assign n659 = g48;
  assign n669 = g4;
  assign n679 = g911;
  assign n684 = g1220;
  assign n689 = g1229;
  assign n694 = g901;
  assign n699 = g2;
  assign n704 = g926;
  assign n709 = g1012;
  assign n719 = g114;
  assign n724 = g134;
  assign n734 = g1524;
  assign n754 = g2;
  assign n759 = g1160;
  assign n774 = g196;
  assign n779 = g48;
  assign n794 = g890;
  assign n804 = g4;
  assign n819 = g1227;
  assign n844 = g48;
  assign n874 = g1284;
  assign n889 = g2;
  assign n894 = g43;
  assign n898 = g8;
  assign n928 = g168;
  assign n938 = g1236;
  assign n943 = g1214;
  assign n953 = g1211;
  assign n958 = g2;
  assign n963 = g110;
  assign n968 = g130;
  assign n973 = g187;
  assign n983 = g1308;
  assign n998 = g8;
  assign n1023 = g1200;
  assign n1027 = g48;
  assign n1042 = g199;
  assign n1052 = g1214;
  assign n1057 = g5;
  assign n1062 = g5;
  assign n1092 = g1270;
  assign n1102 = g906;
  assign n1122 = g1155;
  assign n1132 = g1288;
  assign n1147 = g966;
  assign n1152 = g7;
  assign n1172 = g1207;
  assign n1176 = g906;
  assign n1186 = g2;
  assign n1206 = g1198;
  assign n1211 = g7;
  assign n1231 = ~g1260;
  assign n1236 = g48;
  assign n1246 = g1220;
  assign n1251 = g3;
  assign n1261 = g48;
  assign n1281 = g1206;
  assign n1285 = g1207;
  assign n1290 = g7;
  assign n1295 = g3;
  assign n1300 = g1404;
  assign n1310 = g48;
  assign n1335 = g916;
  assign n1340 = g1424;
  assign n1345 = g1292;
  assign n1355 = g8;
  assign n1374 = g109;
  assign n1379 = g4;
  assign n1403 = g2;
  assign n1408 = g3;
  assign n1418 = g3;
  assign n1438 = g1225;
  assign n1443 = g1250;
  assign n1448 = g138;
  assign n1458 = g48;
  assign n1478 = g1214;
  assign n1483 = g1227;
  assign n1502 = g1196;
  assign n1511 = g28;
  assign n1516 = g530;
  assign n1546 = g7;
  assign n1556 = g45;
  assign n1566 = g1005;
  assign n1585 = g104;
  assign n1590 = g142;
  assign n1595 = g1229;
  assign n1605 = g1224;
  assign n1615 = g1224;
  assign n1645 = g1224;
  assign n1660 = g1227;
  assign n1665 = g1220;
  assign n1669 = g646;
  assign n1679 = g29;
  assign n1689 = g5;
  assign n1699 = g1230;
  assign n1704 = g896;
  assign n1709 = g1225;
  assign n1734 = g6;
  assign n1744 = g4;
  assign n1749 = g891;
  assign n1759 = g1229;
  assign n1764 = g1084;
  assign n1768 = g92;
  assign n1778 = g3;
  assign n1788 = g1234;
  assign n1803 = ~g1252;
  assign n1808 = g1207;
  assign n1822 = g1146;
  assign n1827 = g1229;
  assign n1832 = g95;
  assign n1847 = g1202;
  assign n1851 = g1226;
  assign n1856 = g1217;
  assign n1860 = g1014;
  assign n1895 = g368;
  assign n1930 = g3;
  assign n1945 = g1251;
  assign n1950 = g2;
  assign n1955 = g1081;
  assign n1965 = g1226;
  assign n1980 = g1073;
  assign n2014 = g1156;
  assign n2024 = g1228;
  assign n2029 = g48;
  assign n2034 = g883;
  assign n2044 = g1211;
  assign n2073 = g287;
  assign n2088 = g5;
  assign n2107 = g1403;
  assign n2111 = g89;
  assign n2121 = g1194;
  assign n2140 = g5;
  assign n2145 = g1217;
  assign n2160 = g1228;
  assign n2170 = g5;
  assign n2210 = g1231;
  assign n2215 = g3;
  assign n2225 = g1220;
  assign n2229 = g878;
  assign n2234 = g1198;
  assign n2252 = g1309;
  assign n2257 = g1226;
  assign n2262 = g979;
  assign n2271 = g1240;
  assign n2274 = g891;
  assign n2279 = g48;
  assign n2284 = g1300;
  assign n2289 = g27;
  assign n2298 = g921;
  assign n2313 = g5;
  assign n2318 = g100;
  assign n2328 = g1296;
  assign n2338 = g7;
  assign n2358 = g941;
  assign n2388 = g126;
  assign n2393 = g901;
  assign n2398 = g3;
  assign n2403 = g1191;
  assign n2413 = g26;
  assign n2423 = g94;
  assign n2433 = g1194;
  assign n2438 = g1243;
  assign n2443 = g1260;
  assign n2467 = g1004;
  assign n2475 = g896;
  assign n2478 = g1271;
  assign n2512 = g1226;
  assign n2517 = g4;
  assign n2522 = g7;
  assign n2527 = g1228;
  assign n2532 = g1223;
  assign n2537 = g24;
  assign n2542 = g6236;
  assign n2547 = g6;
  assign n2566 = g1244;
  assign n2581 = g105;
  assign n2586 = g4;
  assign n2591 = g2;
  assign n2610 = g911;
  assign n2619 = g1217;
  assign n2624 = g5;
  assign n2638 = g99;
  assign n2653 = g921;
  assign n2668 = g8;
  assign n2673 = g6;
  assign n2718 = g23;
  assign n2722 = g1393;
  assign n2727 = g1230;
  assign n2732 = g1207;
  assign n2762 = g6;
  assign n2775 = g1185;
  assign n2780 = g1272;
  assign n2784 = g1153;
  assign n2804 = g118;
  assign n2814 = g6;
  assign n2824 = g1311;
  assign n2828 = g4;
  assign n2833 = g207;
  assign n2837 = g1399;
  assign n2847 = g1267;
  assign n2862 = g8;
  assign n2882 = g1223;
  assign n2887 = g1;
  assign n2896 = g1396;
  assign n2901 = g1206;
  assign n2906 = g1224;
  assign n2911 = g7;
  assign n2931 = g122;
  assign n2936 = g202;
  assign n2941 = g37;
  assign n2945 = g576;
  assign n2968 = g1182;
  assign n2982 = g1173;
  assign n2991 = g200;
  assign n3021 = g5;
  assign n3035 = g1199;
  assign n3043 = g1402;
  assign n3052 = g22;
  assign n3055 = g1390;
  assign n3060 = g1034;
  assign n3065 = ~g1260;
  assign n3069 = g1157;
  assign n3089 = g1223;
  assign n3094 = g2;
  assign n3109 = g1214;
  assign n3114 = g1202;
  assign n3124 = g1206;
  assign n3143 = g6;
  assign n3153 = g1240;
  assign n3173 = g8;
  assign n3178 = g2;
  assign n3183 = g1167;
  assign n3202 = g1147;
  assign n3211 = g1154;
  assign n3240 = g3;
  assign n3249 = g1170;
  assign n3268 = g1227;
  assign n3282 = g1192;
  assign n3286 = g16;
  assign n3315 = g1276;
  assign n3329 = g1159;
  assign n3338 = g1310;
  assign n3352 = g4;
  assign n3376 = g3;
  assign n3405 = g1203;
  assign n3449 = g4;
  assign n3464 = g1211;
  assign n3468 = g963;
  assign n3482 = g201;
  assign n3492 = g6;
  assign n3506 = g1163;
  assign n3524 = g1186;
  assign n3534 = g7048;
  assign n3539 = g3;
  always @ (posedge clock) begin
    g397 <= n430;
    g1271 <= n435;
    g312 <= n440;
    g273 <= n445;
    g452 <= n450;
    g948 <= n455;
    g629 <= n460;
    g207 <= n465;
    g1541 <= n470;
    g1153 <= n475;
    g940 <= n480;
    g976 <= n485;
    g498 <= n490;
    g314 <= n495;
    g1092 <= n500;
    g454 <= n505;
    g196 <= n510;
    g535 <= n515;
    g292 <= n520;
    g772 <= n525;
    g1375 <= n530;
    g689 <= n535;
    g183 <= n540;
    g359 <= n545;
    g1384 <= n550;
    g1339 <= n555;
    g20 <= n560;
    g1424 <= n565;
    g767 <= n570;
    g393 <= n575;
    g1077 <= n580;
    g1231 <= n585;
    g294 <= n590;
    g1477 <= n595;
    g4 <= n600;
    g608 <= n605;
    g1205 <= n610;
    g465 <= n614;
    g774 <= n619;
    g921 <= n624;
    g1304 <= n629;
    g243 <= n634;
    g1499 <= n639;
    g80 <= n644;
    g1444 <= n649;
    g1269 <= n654;
    g600 <= n659;
    g423 <= n664;
    g771 <= n669;
    g803 <= n674;
    g843 <= n679;
    g315 <= n684;
    g455 <= n689;
    g906 <= n694;
    g622 <= n699;
    g891 <= n704;
    g1014 <= n709;
    g984 <= n714;
    g117 <= n719;
    g137 <= n724;
    g527 <= n729;
    g1513 <= n734;
    g278 <= n739;
    g1378 <= n744;
    g718 <= n749;
    g598 <= n754;
    g1182 <= n759;
    g1288 <= n764;
    g1382 <= n769;
    g179 <= n774;
    g624 <= n779;
    g48 <= n784;
    g362 <= n789;
    g878 <= n794;
    g270 <= n799;
    g763 <= n804;
    g710 <= n809;
    g730 <= n814;
    g295 <= n819;
    g1037 <= n824;
    g1102 <= n829;
    g483 <= n834;
    g775 <= n839;
    g621 <= n844;
    g1364 <= n849;
    g1454 <= n854;
    g1296 <= n859;
    g5 <= n864;
    g1532 <= n869;
    g587 <= n874;
    g741 <= n879;
    g13 <= n884;
    g606 <= n889;
    g1012 <= n894;
    g52 <= n898;
    g646 <= n903;
    g1412 <= n908;
    g327 <= n913;
    g1189 <= n918;
    g1389 <= n923;
    g1029 <= n928;
    g1371 <= n933;
    g1429 <= n938;
    g398 <= n943;
    g985 <= n948;
    g354 <= n953;
    g619 <= n958;
    g113 <= n963;
    g133 <= n968;
    g180 <= n973;
    g1138 <= n978;
    g1309 <= n983;
    g889 <= n988;
    g390 <= n993;
    g625 <= n998;
    g417 <= n1003;
    g681 <= n1008;
    g437 <= n1013;
    g351 <= n1018;
    g1201 <= n1023;
    g109 <= n1027;
    g1049 <= n1032;
    g1098 <= n1037;
    g200 <= n1042;
    g240 <= n1047;
    g479 <= n1052;
    g126 <= n1057;
    g596 <= n1062;
    g1268 <= n1067;
    g222 <= n1072;
    g420 <= n1077;
    g3 <= n1082;
    g58 <= n1087;
    g172 <= n1092;
    g387 <= n1097;
    g840 <= n1102;
    g365 <= n1107;
    g1486 <= n1112;
    g1504 <= n1117;
    g1185 <= n1122;
    g1385 <= n1127;
    g583 <= n1132;
    g822 <= n1137;
    g1025 <= n1142;
    g969 <= n1147;
    g768 <= n1152;
    g174 <= n1157;
    g685 <= n1162;
    g1087 <= n1167;
    g355 <= n1172;
    g911 <= n1176;
    g1226 <= n1181;
    g99 <= n1186;
    g1045 <= n1191;
    g1173 <= n1196;
    g1373 <= n1201;
    g186 <= n1206;
    g760 <= n1211;
    g959 <= n1216;
    g1369 <= n1221;
    g1007 <= n1226;
    g1459 <= n1231;
    g758 <= n1236;
    g480 <= n1241;
    g396 <= n1246;
    g612 <= n1251;
    g38 <= n1256;
    g632 <= n1261;
    g1415 <= n1266;
    g1227 <= n1271;
    g246 <= n1276;
    g449 <= n1281;
    g517 <= n1285;
    g118 <= n1290;
    g138 <= n1295;
    g16 <= n1300;
    g284 <= n1305;
    g142 <= n1310;
    g219 <= n1315;
    g426 <= n1320;
    g1388 <= n1325;
    g806 <= n1330;
    g846 <= n1335;
    g1428 <= n1340;
    g579 <= n1345;
    g1030 <= n1350;
    g614 <= n1355;
    g1430 <= n1360;
    g1247 <= n1365;
    g669 <= n1370;
    g110 <= n1374;
    g130 <= n1379;
    g225 <= n1384;
    g281 <= n1389;
    g819 <= n1394;
    g1308 <= n1399;
    g611 <= n1403;
    g631 <= n1408;
    g1217 <= n1413;
    g104 <= n1418;
    g1365 <= n1423;
    g825 <= n1428;
    g1333 <= n1433;
    g474 <= n1438;
    g1396 <= n1443;
    g141 <= n1448;
    g1509 <= n1453;
    g766 <= n1458;
    g1018 <= n1463;
    g588 <= n1468;
    g1467 <= n1473;
    g317 <= n1478;
    g457 <= n1483;
    g486 <= n1488;
    g471 <= n1493;
    g1381 <= n1498;
    g1197 <= n1502;
    g513 <= n1506;
    g1397 <= n1511;
    g533 <= n1516;
    g1021 <= n1521;
    g1421 <= n1526;
    g952 <= n1531;
    g1263 <= n1536;
    g580 <= n1541;
    g615 <= n1546;
    g1257 <= n1551;
    g46 <= n1556;
    g402 <= n1561;
    g998 <= n1566;
    g1041 <= n1571;
    g297 <= n1576;
    g954 <= n1581;
    g105 <= n1585;
    g145 <= n1590;
    g212 <= n1595;
    g1368 <= n1600;
    g232 <= n1605;
    g990 <= n1610;
    g475 <= n1615;
    g33 <= n1620;
    g951 <= n1625;
    g799 <= n1630;
    g812 <= n1635;
    g567 <= n1640;
    g313 <= n1645;
    g333 <= n1650;
    g168 <= n1655;
    g214 <= n1660;
    g234 <= n1665;
    g652 <= n1669;
    g1126 <= n1674;
    g1400 <= n1679;
    g1326 <= n1684;
    g92 <= n1689;
    g309 <= n1694;
    g211 <= n1699;
    g834 <= n1704;
    g231 <= n1709;
    g557 <= n1714;
    g1383 <= n1719;
    g1220 <= n1724;
    g158 <= n1729;
    g627 <= n1734;
    g661 <= n1739;
    g77 <= n1744;
    g831 <= n1749;
    g1327 <= n1754;
    g293 <= n1759;
    g1146 <= n1764;
    g89 <= n1768;
    g150 <= n1773;
    g773 <= n1778;
    g859 <= n1783;
    g1240 <= n1788;
    g518 <= n1793;
    g1472 <= n1798;
    g1443 <= n1803;
    g436 <= n1808;
    g405 <= n1813;
    g1034 <= n1818;
    g1147 <= n1822;
    g374 <= n1827;
    g98 <= n1832;
    g563 <= n1837;
    g510 <= n1842;
    g530 <= n1847;
    g215 <= n1851;
    g235 <= n1856;
    g1013 <= n1860;
    g6 <= n1865;
    g55 <= n1870;
    g1317 <= n1875;
    g504 <= n1880;
    g665 <= n1885;
    g544 <= n1890;
    g371 <= n1895;
    g62 <= n1900;
    g792 <= n1905;
    g468 <= n1910;
    g815 <= n1915;
    g1460 <= n1920;
    g553 <= n1925;
    g623 <= n1930;
    g501 <= n1935;
    g1190 <= n1940;
    g1390 <= n1945;
    g74 <= n1950;
    g1156 <= n1955;
    g318 <= n1960;
    g458 <= n1965;
    g342 <= n1970;
    g1250 <= n1975;
    g1163 <= n1980;
    g1363 <= n1985;
    g1432 <= n1990;
    g1053 <= n1995;
    g252 <= n2000;
    g330 <= n2005;
    g264 <= n2010;
    g1157 <= n2014;
    g1357 <= n2019;
    g375 <= n2024;
    g68 <= n2029;
    g852 <= n2034;
    g261 <= n2039;
    g516 <= n2044;
    g536 <= n2049;
    g979 <= n2054;
    g778 <= n2059;
    g199 <= n2064;
    g1292 <= n2068;
    g290 <= n2073;
    g1084 <= n2078;
    g1439 <= n2083;
    g770 <= n2088;
    g1276 <= n2093;
    g890 <= n2098;
    g1004 <= n2102;
    g1404 <= n2107;
    g93 <= n2111;
    g2 <= n2116;
    g287 <= n2121;
    g560 <= n2125;
    g1224 <= n2130;
    g1320 <= n2135;
    g617 <= n2140;
    g316 <= n2145;
    g336 <= n2150;
    g933 <= n2155;
    g456 <= n2160;
    g345 <= n2165;
    g628 <= n2170;
    g8 <= n2175;
    g887 <= n2180;
    g789 <= n2185;
    g173 <= n2190;
    g550 <= n2195;
    g255 <= n2200;
    g949 <= n2205;
    g1244 <= n2210;
    g620 <= n2215;
    g1435 <= n2220;
    g477 <= n2225;
    g926 <= n2229;
    g368 <= n2234;
    g855 <= n2238;
    g1214 <= n2243;
    g1110 <= n2248;
    g1310 <= n2252;
    g296 <= n2257;
    g972 <= n2262;
    g1402 <= n2267;
    g1236 <= n2271;
    g896 <= n2274;
    g613 <= n2279;
    g566 <= n2284;
    g1394 <= n2289;
    g1489 <= n2294;
    g883 <= n2298;
    g47 <= n2303;
    g971 <= n2308;
    g609 <= n2313;
    g103 <= n2318;
    g1254 <= n2323;
    g556 <= n2328;
    g1409 <= n2333;
    g626 <= n2338;
    g1229 <= n2343;
    g782 <= n2348;
    g237 <= n2353;
    g942 <= n2358;
    g228 <= n2363;
    g706 <= n2368;
    g746 <= n2373;
    g1462 <= n2378;
    g963 <= n2383;
    g129 <= n2388;
    g837 <= n2393;
    g599 <= n2398;
    g1192 <= n2403;
    g828 <= n2408;
    g1392 <= n2413;
    g492 <= n2418;
    g95 <= n2423;
    g944 <= n2428;
    g195 <= n2433;
    g1431 <= n2438;
    g1252 <= n2443;
    g356 <= n2448;
    g953 <= n2453;
    g1176 <= n2458;
    g1376 <= n2463;
    g1005 <= n2467;
    g1405 <= n2471;
    g901 <= n2475;
    g1270 <= n2478;
    g1225 <= n2482;
    g1073 <= n2487;
    g1324 <= n2492;
    g1069 <= n2497;
    g443 <= n2502;
    g1377 <= n2507;
    g377 <= n2512;
    g618 <= n2517;
    g602 <= n2522;
    g213 <= n2527;
    g233 <= n2532;
    g1199 <= n2537;
    g1399 <= n2542;
    g83 <= n2547;
    g888 <= n2552;
    g573 <= n2557;
    g399 <= n2562;
    g1245 <= n2566;
    g507 <= n2571;
    g547 <= n2576;
    g108 <= n2581;
    g610 <= n2586;
    g630 <= n2591;
    g1207 <= n2596;
    g249 <= n2601;
    g65 <= n2606;
    g916 <= n2610;
    g936 <= n2614;
    g478 <= n2619;
    g604 <= n2624;
    g945 <= n2629;
    g1114 <= n2634;
    g100 <= n2638;
    g429 <= n2643;
    g809 <= n2648;
    g849 <= n2653;
    g1408 <= n2658;
    g1336 <= n2663;
    g601 <= n2668;
    g122 <= n2673;
    g1065 <= n2678;
    g1122 <= n2683;
    g1228 <= n2688;
    g495 <= n2693;
    g1322 <= n2698;
    g1230 <= n2703;
    g1033 <= n2708;
    g267 <= n2713;
    g1195 <= n2718;
    g1395 <= n2722;
    g373 <= n2727;
    g274 <= n2732;
    g1266 <= n2737;
    g714 <= n2742;
    g734 <= n2747;
    g1142 <= n2752;
    g1342 <= n2757;
    g769 <= n2762;
    g1081 <= n2767;
    g1481 <= n2771;
    g1097 <= n2775;
    g543 <= n2780;
    g1154 <= n2784;
    g1354 <= n2789;
    g489 <= n2794;
    g874 <= n2799;
    g121 <= n2804;
    g591 <= n2809;
    g616 <= n2814;
    g1267 <= n2819;
    g1312 <= n2824;
    g605 <= n2828;
    g182 <= n2833;
    g1401 <= n2837;
    g950 <= n2842;
    g1329 <= n2847;
    g408 <= n2852;
    g871 <= n2857;
    g759 <= n2862;
    g146 <= n2867;
    g202 <= n2872;
    g440 <= n2877;
    g476 <= n2882;
    g184 <= n2887;
    g1149 <= n2892;
    g1398 <= n2896;
    g210 <= n2901;
    g394 <= n2906;
    g86 <= n2911;
    g570 <= n2916;
    g275 <= n2921;
    g303 <= n2926;
    g125 <= n2931;
    g181 <= n2936;
    g1524 <= n2941;
    g595 <= n2945;
    g1319 <= n2950;
    g863 <= n2955;
    g1211 <= n2960;
    g966 <= n2965;
    g1186 <= n2968;
    g1386 <= n2973;
    g875 <= n2978;
    g1170 <= n2982;
    g1370 <= n2987;
    g201 <= n2991;
    g1325 <= n2996;
    g1280 <= n3001;
    g1106 <= n3006;
    g1061 <= n3011;
    g1387 <= n3016;
    g762 <= n3021;
    g1461 <= n3026;
    g378 <= n3031;
    g1200 <= n3035;
    g1514 <= n3039;
    g1403 <= n3043;
    g1345 <= n3047;
    g1191 <= n3052;
    g1391 <= n3055;
    g185 <= n3060;
    g1307 <= n3065;
    g1159 <= n3069;
    g1223 <= n3074;
    g446 <= n3079;
    g1416 <= n3084;
    g395 <= n3089;
    g764 <= n3094;
    g1251 <= n3099;
    g216 <= n3104;
    g236 <= n3109;
    g205 <= n3114;
    g540 <= n3119;
    g576 <= n3124;
    g1537 <= n3128;
    g727 <= n3133;
    g999 <= n3138;
    g761 <= n3143;
    g1272 <= n3148;
    g1243 <= n3153;
    g1328 <= n3158;
    g1130 <= n3163;
    g1330 <= n3168;
    g114 <= n3173;
    g134 <= n3178;
    g1166 <= n3183;
    g524 <= n3188;
    g1366 <= n3193;
    g348 <= n3198;
    g1148 <= n3202;
    g1348 <= n3207;
    g1155 <= n3211;
    g1260 <= n3215;
    g7 <= n3220;
    g258 <= n3225;
    g521 <= n3230;
    g300 <= n3235;
    g765 <= n3240;
    g1118 <= n3245;
    g1167 <= n3249;
    g1318 <= n3253;
    g1367 <= n3258;
    g677 <= n3263;
    g376 <= n3268;
    g1057 <= n3273;
    g973 <= n3278;
    g1193 <= n3282;
    g1393 <= n3286;
    g1549 <= n3290;
    g1321 <= n3295;
    g1253 <= n3300;
    g1519 <= n3305;
    g584 <= n3310;
    g539 <= n3315;
    g324 <= n3320;
    g432 <= n3325;
    g1158 <= n3329;
    g321 <= n3334;
    g1311 <= n3338;
    g414 <= n3342;
    g1374 <= n3347;
    g94 <= n3352;
    g1284 <= n3356;
    g1545 <= n3361;
    g1380 <= n3366;
    g673 <= n3371;
    g607 <= n3376;
    g306 <= n3381;
    g943 <= n3386;
    g162 <= n3391;
    g411 <= n3396;
    g866 <= n3401;
    g1204 <= n3405;
    g1300 <= n3409;
    g384 <= n3414;
    g339 <= n3419;
    g459 <= n3424;
    g1323 <= n3429;
    g381 <= n3434;
    g1528 <= n3439;
    g1351 <= n3444;
    g597 <= n3449;
    g1372 <= n3454;
    g154 <= n3459;
    g435 <= n3464;
    g970 <= n3468;
    g1134 <= n3473;
    g995 <= n3478;
    g190 <= n3482;
    g1313 <= n3487;
    g603 <= n3492;
    g1494 <= n3497;
    g462 <= n3502;
    g1160 <= n3506;
    g1360 <= n3510;
    g1450 <= n3515;
    g187 <= n3520;
    g1179 <= n3524;
    g1379 <= n3529;
    g12 <= n3534;
    g71 <= n3539;
  end
endmodule


