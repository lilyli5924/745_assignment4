module medium_2 ( clock, 
    g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558,
    g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39,
    g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23,
    g2584, g3222, g3600, g4307, g4321, g4422, g4809, g5137, g5468, g5469,
    g5692, g6282, g6284, g6360, g6362, g6364, g6366, g6368, g6370, g6372,
    g6374, g6728, g1290, g4121, g4108, g4106, g4103, g1293, g4099, g4102,
    g4109, g4100, g4112, g4105, g4101, g4110, g4104, g4107, g4098  );
  input  clock, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557,
    g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42,
    g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23;
  output g2584, g3222, g3600, g4307, g4321, g4422, g4809, g5137, g5468, g5469,
    g5692, g6282, g6284, g6360, g6362, g6364, g6366, g6368, g6370, g6372,
    g6374, g6728, g1290, g4121, g4108, g4106, g4103, g1293, g4099, g4102,
    g4109, g4100, g4112, g4105, g4101, g4110, g4104, g4107, g4098;
  reg g678, g332, g123, g207, g695, g461, g18, g292, g331, g689, g24, g465,
    g84, g291, g676, g622, g117, g278, g128, g598, g554, g496, g179, g48,
    g590, g551, g682, g11, g606, g188, g646, g327, g361, g289, g398, g684,
    g619, g208, g248, g390, g625, g681, g437, g276, g3, g323, g224, g685,
    g43, g157, g282, g697, g206, g449, g118, g528, g284, g426, g634, g669,
    g520, g281, g175, g15, g631, g69, g693, g337, g457, g486, g471, g328,
    g285, g418, g402, g297, g212, g410, g430, g33, g662, g453, g269, g574,
    g441, g664, g349, g211, g586, g571, g29, g326, g698, g654, g293, g690,
    g445, g374, g6, g687, g357, g386, g504, g665, g166, g541, g74, g338,
    g696, g516, g536, g683, g353, g545, g254, g341, g290, g2, g287, g336,
    g345, g628, g679, g28, g688, g283, g613, g10, g14, g680, g143, g672,
    g667, g366, g279, g492, g170, g686, g288, g638, g602, g642, g280, g663,
    g610, g148, g209, g675, g478, g122, g54, g594, g286, g489, g616, g79,
    g218, g242, g578, g184, g119, g668, g139, g422, g210, g394, g230, g25,
    g204, g658, g650, g378, g508, g548, g370, g406, g236, g500, g205, g197,
    g666, g114, g524, g260, g111, g131, g7, g19, g677, g582, g485, g699,
    g193, g135, g382, g414, g434, g266, g49, g152, g692, g277, g127, g161,
    g512, g532, g64, g694, g691, g1, g59;
  wire n711_1, n712, n713, n714, n715, n716_1, n717, n718, n719, n720,
    n721_1, n722, n723, n724, n725, n726_1, n727, n728, n729, n730, n731_1,
    n732, n733, n734, n735, n736_1, n737, n738, n739, n741_1, n742, n743,
    n744, n745, n746_1, n747, n748, n749, n750, n751_1, n752, n753, n754,
    n755, n756_1, n757, n758, n759, n760, n761_1, n762, n763, n773, n775,
    n776_1, n777, n778, n779, n780, n781_1, n782, n783, n784, n785, n786_1,
    n787, n788, n789, n790, n791_1, n792, n793, n794, n795, n796_1, n797,
    n798, n799, n800, n801_1, n802, n803, n805, n806_1, n807, n808, n809,
    n810, n811_1, n812, n813, n814, n815, n816_1, n817, n818, n819, n820,
    n821_1, n822, n823, n824, n825, n826_1, n827, n828, n829, n830, n831_1,
    n832, n833, n834, n835, n836_1, n837, n838, n839, n840, n841_1, n842,
    n843, n844, n845, n846_1, n847, n848, n849, n850, n851_1, n852, n853,
    n854, n855, n856_1, n857, n858, n859, n860, n861_1, n862, n863, n864,
    n865, n866_1, n867, n868, n869, n870, n871_1, n872, n873, n874, n875,
    n876_1, n877, n878, n879, n880, n881_1, n882, n883, n884, n885, n886_1,
    n887, n888, n889, n890, n891_1, n892, n893, n894, n895, n896_1, n897,
    n898, n899, n900, n901_1, n902, n903, n904, n905, n906_1, n907, n908,
    n909, n910, n911_1, n912, n913, n914, n915, n916_1, n917, n918, n919,
    n920, n921_1, n922, n923, n924, n925, n926_1, n927, n928, n929, n930,
    n931_1, n932, n933, n934, n935, n936_1, n937, n938, n939, n940, n941_1,
    n942, n943, n944, n945, n946_1, n947, n948, n949, n950, n951_1, n952,
    n953, n954, n955, n956_1, n957, n958, n959, n960, n961_1, n962, n963,
    n964, n965, n966_1, n967, n968, n969, n970, n971_1, n972, n973, n974,
    n975, n976_1, n977, n978, n979, n980, n981_1, n982, n983, n984, n986_1,
    n987, n988, n989, n990, n991_1, n992, n993, n994, n995, n996_1, n997,
    n998, n999, n1000, n1001_1, n1002, n1003, n1004, n1005, n1006_1, n1007,
    n1008, n1009, n1010, n1011_1, n1012, n1013, n1014, n1015, n1016_1,
    n1018, n1019, n1021_1, n1022, n1023, n1024, n1025, n1027, n1028, n1029,
    n1030, n1031_1, n1032, n1033, n1034, n1035, n1036_1, n1037, n1038,
    n1039, n1040, n1041_1, n1042, n1043, n1044, n1045, n1046_1, n1047,
    n1048, n1049, n1050, n1051_1, n1052, n1053, n1054, n1055, n1056_1,
    n1057, n1058, n1059, n1060, n1061_1, n1062, n1063, n1064, n1065,
    n1066_1, n1067, n1068, n1069, n1070, n1071_1, n1072, n1073, n1074,
    n1075, n1076_1, n1077, n1079, n1080, n1081_1, n1082, n1083, n1084,
    n1086_1, n1087, n1088, n1089, n1090, n1091_1, n1092, n1093, n1094,
    n1095, n1097, n1098, n1099, n1101_1, n1102, n1103, n1105, n1106_1,
    n1108, n1109, n1110, n1111_1, n1112, n1113, n1114, n1115, n1116_1,
    n1117, n1118, n1119, n1120, n1121_1, n1122, n1123, n1124, n1125,
    n1126_1, n1127, n1128, n1129, n1130, n1131_1, n1132, n1133, n1134,
    n1136_1, n1137, n1138, n1139, n1140, n1141_1, n1142, n1143, n1144,
    n1145, n1146_1, n1147, n1148, n1149, n1150, n1151_1, n1152, n1153,
    n1154, n1155, n1156_1, n1157, n1158, n1159, n1160, n1161_1, n1162,
    n1163, n1164, n1165, n1166_1, n1168, n1169, n1170, n1171_1, n1172,
    n1173, n1174, n1175, n1176_1, n1177, n1178, n1179, n1181_1, n1182,
    n1184, n1185, n1186_1, n1187, n1188, n1189, n1190, n1191_1, n1192,
    n1193, n1194, n1195, n1196_1, n1197, n1198, n1199, n1200, n1201_1,
    n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
    n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1228, n1229, n1230, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1240, n1241, n1244, n1245, n1246,
    n1247, n1248, n1249, n1251, n1252, n1253, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1264, n1265, n1267, n1269, n1270, n1271,
    n1272, n1273, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1317, n1318, n1319, n1320, n1321, n1322, n1324, n1325, n1328,
    n1329, n1330, n1332, n1333, n1335, n1337, n1339, n1340, n1341, n1342,
    n1343, n1344, n1345, n1346, n1347, n1348, n1350, n1351, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1375,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1388,
    n1389, n1392, n1393, n1395, n1396, n1397, n1398, n1399, n1401, n1402,
    n1403, n1405, n1406, n1408, n1409, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1441, n1442, n1444, n1445, n1447, n1448,
    n1450, n1451, n1453, n1454, n1455, n1456, n1458, n1460, n1461, n1462,
    n1463, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1484, n1486,
    n1487, n1489, n1490, n1492, n1493, n1495, n1496, n1498, n1499, n1501,
    n1502, n1504, n1505, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
    n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1525,
    n1526, n1528, n1529, n1531, n1532, n1533, n1534, n1535, n1537, n1538,
    n1540, n1541, n1543, n1544, n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
    n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
    n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
    n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
    n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
    n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1662,
    n1663, n1665, n1667, n1668, n1670, n1671, n1672, n1673, n1674, n1675,
    n1677, n1679, n1680, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1702,
    n1703, n1704, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
    n1727, n1729, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
    n1739, n1741, n1743, n1744, n1746, n1748, n1749, n1751, n1752, n1754,
    n1755, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
    n1766, n1767, n1768, n1771, n1773, n1774, n1776, n1777, n1779, n1780,
    n1782, n1783, n1785, n1786, n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1797, n1798, n1801, n1802, n1804, n1805, n1806, n1808,
    n1809, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
    n1830, n1831, n1832, n1833, n1834, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1849, n1851, n1852,
    n1854, n1855, n1857, n1858, n1860, n1861, n1863, n1864, n1867, n1868,
    n1869, n1870, n1871, n1872, n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1917, n1918, n1920, n1921, n1923, n1924,
    n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941, n151, n156, n161, n166, n171,
    n176, n181, n186, n191, n196, n201, n206, n211, n216, n221, n226, n231,
    n236, n241, n246, n251, n256, n261, n266, n271, n276, n281, n286, n291,
    n296, n301, n306, n311, n316, n321, n326, n331, n336, n341, n346, n351,
    n356, n361, n366, n371, n376, n381, n386, n391, n396, n401, n406, n411,
    n416, n421, n426, n431, n436, n441, n446, n451, n456, n461, n466, n471,
    n476, n481, n486, n491, n496, n501, n506, n511, n516, n521, n526, n531,
    n536, n541, n546, n551, n556, n561, n566, n571, n576, n581, n586, n591,
    n596, n601, n606, n611, n616, n621, n626, n631, n636, n641, n646, n651,
    n656, n661, n666, n671, n676, n681, n686, n691, n696, n701, n706, n711,
    n716, n721, n726, n731, n736, n741, n746, n751, n756, n761, n766, n771,
    n776, n781, n786, n791, n796, n801, n806, n811, n816, n821, n826, n831,
    n836, n841, n846, n851, n856, n861, n866, n871, n876, n881, n886, n891,
    n896, n901, n906, n911, n916, n921, n926, n931, n936, n941, n946, n951,
    n956, n961, n966, n971, n976, n981, n986, n991, n996, n1001, n1006,
    n1011, n1016, n1021, n1026, n1031, n1036, n1041, n1046, n1051, n1056,
    n1061, n1066, n1071, n1076, n1081, n1086, n1091, n1096, n1101, n1106,
    n1111, n1116, n1121, n1126, n1131, n1136, n1141, n1146, n1151, n1156,
    n1161, n1166, n1171, n1176, n1181, n1186, n1191, n1196, n1201;
  assign g2584 = g89 & ~g102;
  assign g4809 = ~n711_1 & ~n712;
  assign n711_1 = g496 & ~g486;
  assign n712 = g492 & ~g489;
  assign n713 = ~g22 & g675 & g676 & ~n714;
  assign n714 = ~g41 & ~n715;
  assign n715 = ~n716_1 & ~n739;
  assign n716_1 = g48 & n717;
  assign n717 = ~n718 & ~n738;
  assign n718 = n719 & ~n725;
  assign n719 = ~n720 & ~n724;
  assign n720 = g18 & ~n721_1;
  assign n721_1 = ~n722 & ~n723;
  assign n722 = g24 & ~g28;
  assign n723 = ~g24 & g28;
  assign n724 = ~g18 & n721_1;
  assign n725 = ~n726_1 & ~n737;
  assign n726_1 = g14 & ~n727;
  assign n727 = ~n728 & ~n736_1;
  assign n728 = n729 & n733;
  assign n729 = ~n730 & ~n732;
  assign n730 = g1 & ~n731_1;
  assign n731_1 = g2 & g1;
  assign n732 = g2 & ~n731_1;
  assign n733 = ~n734 & ~n735;
  assign n734 = g6 & ~g10;
  assign n735 = ~g6 & g10;
  assign n736_1 = ~n729 & ~n733;
  assign n737 = ~g14 & n727;
  assign n738 = ~n719 & n725;
  assign n739 = ~g48 & ~n717;
  assign g6284 = ~n741_1 | ~n742;
  assign n741_1 = g41 & n713;
  assign n742 = ~n743 & ~n763;
  assign n743 = n744 & ~n750;
  assign n744 = ~n745 & ~n749;
  assign n745 = g11 & ~n746_1;
  assign n746_1 = ~n747 & ~n748;
  assign n747 = g3 & ~g7;
  assign n748 = ~g3 & g7;
  assign n749 = ~g11 & n746_1;
  assign n750 = ~n751_1 & ~n762;
  assign n751_1 = g15 & ~n752;
  assign n752 = ~n753 & ~n761_1;
  assign n753 = n754 & n758;
  assign n754 = ~n755 & ~n757;
  assign n755 = g33 & ~n756_1;
  assign n756_1 = g33 & g29;
  assign n757 = g29 & ~n756_1;
  assign n758 = ~n759 & ~n760;
  assign n759 = g25 & ~g19;
  assign n760 = ~g25 & g19;
  assign n761_1 = ~n754 & ~n758;
  assign n762 = ~g15 & n752;
  assign n763 = ~n744 & n750;
  assign g6360 = g25 | ~n741_1;
  assign g6362 = g29 | ~n741_1;
  assign g6364 = g3 | ~n741_1;
  assign g6366 = g33 | ~n741_1;
  assign g6368 = g7 | ~n741_1;
  assign g6370 = g11 | ~n741_1;
  assign g6372 = g15 | ~n741_1;
  assign g6374 = g19 | ~n741_1;
  assign g4121 = ~g638 | n773;
  assign n773 = ~g567 & g638;
  assign n156 = n775 | n788;
  assign n775 = ~n776_1 & ~n777 & ~n781_1;
  assign n776_1 = ~g314 & ~g301 & ~g310 & ~g306;
  assign n777 = g332 & n778;
  assign n778 = g323 & ~g357 & n779;
  assign n779 = ~g353 & ~g349 & n780;
  assign n780 = ~g345 & ~g338 & ~g341;
  assign n781_1 = ~g332 & ~n782;
  assign n782 = n778 & ~n783;
  assign n783 = ~n787 & ~n784 & ~n785 & ~n786_1;
  assign n784 = g310 & g314;
  assign n785 = g306 & ~g310;
  assign n786_1 = g306 & ~g314;
  assign n787 = ~g306 & g310 & ~g314;
  assign n788 = n776_1 & ~n789;
  assign n789 = ~g337 & ~n790 & ~n800;
  assign n790 = ~n791_1 & ~n792 & ~n796_1;
  assign n791_1 = g662 & g658;
  assign n792 = ~g687 & n793 & n795;
  assign n793 = ~n714 & g676 & n794 & g41 & g702 & g699;
  assign n794 = g662 & ~g658;
  assign n795 = g689 & ~g698;
  assign n796_1 = n795 & n797;
  assign n797 = ~g687 & n798;
  assign n798 = n794 & n799;
  assign n799 = g699 & g702 & ~g41 & g676 & ~n714;
  assign n800 = ~n791_1 & ~n801_1 & ~n802;
  assign n801_1 = n795 & g687 & n793;
  assign n802 = n795 & n803;
  assign n803 = g687 & n798;
  assign n161 = n805 | n817;
  assign n805 = ~n806_1 & ~n807 & ~n810;
  assign n806_1 = ~g102 & ~g89 & ~g98 & ~g94;
  assign n807 = g123 & n808;
  assign n808 = g114 & ~g139 & n809;
  assign n809 = ~g135 & ~g128 & ~g131;
  assign n810 = ~g123 & ~n811_1;
  assign n811_1 = n808 & ~n812;
  assign n812 = ~n816_1 & ~n813 & ~n814 & ~n815;
  assign n813 = g98 & g102;
  assign n814 = g94 & ~g98;
  assign n815 = g94 & ~g102;
  assign n816_1 = ~g94 & g98 & ~g102;
  assign n817 = n806_1 & ~n818;
  assign n818 = ~n841_1 & ~n819 & ~n823 & ~n838;
  assign n819 = ~n791_1 & ~n820 & ~n822;
  assign n820 = n793 & ~g685 & n821_1 & g684;
  assign n821_1 = ~g688 & g689 & g698;
  assign n822 = n798 & n821_1 & ~g685 & g684;
  assign n823 = ~n824 & ~n831_1;
  assign n824 = ~n825 & ~n828;
  assign n825 = ~n826_1 & ~n827;
  assign n826_1 = g658 & g650;
  assign n827 = g681 & ~g658;
  assign n828 = ~n829 & ~n830;
  assign n829 = g646 & g658;
  assign n830 = g680 & ~g658;
  assign n831_1 = ~n832 & ~n835;
  assign n832 = ~n833 & ~n834;
  assign n833 = g606 & g658;
  assign n834 = g679 & ~g658;
  assign n835 = ~n836_1 & ~n837;
  assign n836_1 = g642 & g658;
  assign n837 = g678 & ~g658;
  assign n838 = ~n839 & ~n840;
  assign n839 = g658 & g260;
  assign n840 = g686 & ~g658;
  assign n841_1 = ~n842 & ~n862 & ~n963;
  assign n842 = ~n843 & ~n858;
  assign n843 = ~n844 & ~n851_1;
  assign n844 = ~n845 & ~n848;
  assign n845 = ~n846_1 & ~n847;
  assign n846_1 = g254 & g658;
  assign n847 = g685 & ~g658;
  assign n848 = ~n849 & ~n850;
  assign n849 = g248 & g658;
  assign n850 = g684 & ~g658;
  assign n851_1 = ~n852 & ~n855;
  assign n852 = ~n853 & ~n854;
  assign n853 = g683 & ~g658;
  assign n854 = g242 & g658;
  assign n855 = ~n856_1 & ~n857;
  assign n856_1 = g682 & ~g658;
  assign n857 = g658 & g236;
  assign n858 = ~n859 & ~n860;
  assign n859 = g297 & n791_1;
  assign n860 = n803 & n861_1 & g688;
  assign n861_1 = ~g689 & ~g698;
  assign n862 = g658 & ~n863;
  assign n863 = ~n864 & n910;
  assign n864 = ~n865 & ~n882;
  assign n865 = ~n880 & ~n874 & ~n866_1 & ~n867 & ~n872 & ~n875;
  assign n866_1 = g692 & ~g567 & g598 & ~g634;
  assign n867 = ~g598 & ~n868 & ~n870;
  assign n868 = ~g567 & ~n869;
  assign n869 = ~g634 & g690;
  assign n870 = g567 & ~n871_1;
  assign n871_1 = ~g634 & g691;
  assign n872 = ~g634 & g693 & n873;
  assign n873 = g567 & g598;
  assign n874 = ~g567 & g598 & g634 & g696;
  assign n875 = ~g598 & ~n876_1 & ~n878;
  assign n876_1 = ~g567 & ~n877;
  assign n877 = g634 & g694;
  assign n878 = g567 & ~n879;
  assign n879 = g695 & g634;
  assign n880 = g697 & n881_1;
  assign n881_1 = g634 & n873;
  assign n882 = ~n898 & ~n892 & ~n883 & ~n886_1 & ~n889 & ~n895 & ~n901_1 & ~n904 & ~n907;
  assign n883 = ~n884 & ~n885;
  assign n884 = g292 & g686;
  assign n885 = ~g292 & ~g686;
  assign n886_1 = ~n887 & ~n888;
  assign n887 = g291 & g685;
  assign n888 = ~g291 & ~g685;
  assign n889 = ~n890 & ~n891_1;
  assign n890 = g684 & g290;
  assign n891_1 = ~g684 & ~g290;
  assign n892 = ~n893 & ~n894;
  assign n893 = g682 & g288;
  assign n894 = ~g682 & ~g288;
  assign n895 = ~n896_1 & ~n897;
  assign n896_1 = g289 & g683;
  assign n897 = ~g289 & ~g683;
  assign n898 = ~n899 & ~n900;
  assign n899 = g681 & g287;
  assign n900 = ~g681 & ~g287;
  assign n901_1 = ~n902 & ~n903;
  assign n902 = g680 & g286;
  assign n903 = ~g680 & ~g286;
  assign n904 = ~n905 & ~n906_1;
  assign n905 = g285 & g679;
  assign n906_1 = ~g285 & ~g679;
  assign n907 = ~n908 & ~n909;
  assign n908 = g678 & g284;
  assign n909 = ~g678 & ~g284;
  assign n910 = ~n911_1 & ~n961_1;
  assign n911_1 = ~n960 & ~n912 & ~n958 & ~n959;
  assign n912 = n928 & ~n913 & ~n922 & g283;
  assign n913 = ~g282 & ~g283 & n914;
  assign n914 = ~g478 & n915;
  assign n915 = ~n916_1 & ~n920;
  assign n916_1 = ~n917 & ~n919;
  assign n917 = g281 & ~n918;
  assign n918 = g281 & g280;
  assign n919 = g280 & ~n918;
  assign n920 = ~g280 & g281 & n921_1 & g279;
  assign n921_1 = g277 & g276 & g278;
  assign n922 = n923 & n927;
  assign n923 = ~n916_1 & ~n924;
  assign n924 = ~n914 & ~n925;
  assign n925 = g478 & ~n926_1;
  assign n926_1 = g478 & n915;
  assign n927 = g282 & ~g283;
  assign n928 = ~n955 & ~n929 & ~n931_1 & ~n932;
  assign n929 = n930 & ~g282 & g283;
  assign n930 = n918 & n921_1 & g279;
  assign n931_1 = ~n915 & ~g282 & ~g283 & ~g478;
  assign n932 = n930 & n933;
  assign n933 = n927 & n934;
  assign n934 = n916_1 & ~n935;
  assign n935 = ~n936_1 & ~n954;
  assign n936_1 = g478 & ~n937;
  assign n937 = ~n938 & ~n946_1;
  assign n938 = g278 & ~n939;
  assign n939 = ~n940 & ~n943;
  assign n940 = ~g277 & ~n941_1 & ~n942;
  assign n941_1 = ~g276 & g693;
  assign n942 = g276 & g692;
  assign n943 = g277 & ~n944 & ~n945;
  assign n944 = ~g276 & g691;
  assign n945 = g276 & g690;
  assign n946_1 = ~g278 & ~n947;
  assign n947 = ~n948 & ~n951_1;
  assign n948 = ~g277 & ~n949 & ~n950;
  assign n949 = ~g276 & g697;
  assign n950 = g276 & g696;
  assign n951_1 = g277 & ~n952 & ~n953;
  assign n952 = g695 & ~g276;
  assign n953 = g276 & g694;
  assign n954 = ~g478 & n937;
  assign n955 = n930 & n956_1;
  assign n956_1 = ~n957 & g282 & g283;
  assign n957 = ~n923 & ~n934;
  assign n958 = ~n930 & n956_1;
  assign n959 = ~n930 & n933;
  assign n960 = ~n933 & n927 & n930;
  assign n961_1 = ~n962 & n928 & ~n960;
  assign n962 = ~n959 & ~n958 & ~n913 & ~n922 & g282;
  assign n963 = g690 & ~g658;
  assign n964 = ~n965 & ~n984;
  assign n965 = g197 & ~n966_1 & ~n974;
  assign n966_1 = ~g210 & ~g471 & ~n967 & ~g211;
  assign n967 = ~n968 & ~n970;
  assign n968 = n969 & g207 & ~g208 & g209;
  assign n969 = g205 & g204 & g206;
  assign n970 = ~n971_1 & ~n973;
  assign n971_1 = g209 & ~n972;
  assign n972 = g208 & g209;
  assign n973 = g208 & ~n972;
  assign n974 = n975 & ~n979;
  assign n975 = ~n976_1 & ~n977;
  assign n976_1 = n972 & n969 & g207;
  assign n977 = ~g211 & ~g210 & n978;
  assign n978 = ~g471 & n967;
  assign n979 = ~n980 & ~n983;
  assign n980 = g207 & n981_1;
  assign n981_1 = g206 & n982;
  assign n982 = g204 & g205;
  assign n983 = ~g207 & ~n981_1;
  assign n984 = g693 & ~g197;
  assign n176 = n986_1 | n1016_1;
  assign n986_1 = g461 & ~n987;
  assign n987 = ~g541 & ~g536 & n988;
  assign n988 = ~n1004 & ~n998 & ~n989 & ~n992 & ~n995 & ~n1001_1 & ~n1007 & ~n1010 & ~n1013;
  assign n989 = ~n990 & ~n991_1;
  assign n990 = g212 & g500;
  assign n991_1 = ~g212 & ~g500;
  assign n992 = ~n993 & ~n994;
  assign n993 = g504 & g218;
  assign n994 = ~g504 & ~g218;
  assign n995 = ~n996_1 & ~n997;
  assign n996_1 = g224 & g508;
  assign n997 = ~g224 & ~g508;
  assign n998 = ~n999 & ~n1000;
  assign n999 = g230 & g512;
  assign n1000 = ~g230 & ~g512;
  assign n1001_1 = ~n1002 & ~n1003;
  assign n1002 = g516 & g236;
  assign n1003 = ~g516 & ~g236;
  assign n1004 = ~n1005 & ~n1006_1;
  assign n1005 = g520 & g242;
  assign n1006_1 = ~g520 & ~g242;
  assign n1007 = ~n1008 & ~n1009;
  assign n1008 = g248 & g524;
  assign n1009 = ~g248 & ~g524;
  assign n1010 = ~n1011_1 & ~n1012;
  assign n1011_1 = g528 & g254;
  assign n1012 = ~g528 & ~g254;
  assign n1013 = ~n1014 & ~n1015;
  assign n1014 = g260 & g532;
  assign n1015 = ~g260 & ~g532;
  assign n1016_1 = g430 & n987;
  assign n191 = g328 & ~n1018;
  assign n1018 = n783 & ~n1019;
  assign n1019 = ~g306 & g314;
  assign n206 = n1021_1 | n1025;
  assign n1021_1 = g465 & ~n1022;
  assign n1022 = ~g677 & n1023;
  assign n1023 = g683 & g684 & n799 & n1024 & ~g682 & ~g681;
  assign n1024 = g685 & n821_1;
  assign n1025 = g691 & n1022;
  assign n211 = n1027 | n1055;
  assign n1027 = n1028 & ~n1044 & ~n1054;
  assign n1028 = ~n776_1 & ~n1029;
  assign n1029 = ~n1030 & ~n1035;
  assign n1030 = ~n1031_1 & ~n1033;
  assign n1031_1 = n777 & ~n1032;
  assign n1032 = ~g306 & ~g310;
  assign n1033 = n778 & n1034;
  assign n1034 = ~g319 & g301 & g314;
  assign n1035 = ~n1036_1 & ~n1041_1;
  assign n1036_1 = ~g84 & n1037;
  assign n1037 = n1039 & ~g54 & ~g64 & ~g79 & ~g74 & ~g69 & ~g59 & n1038;
  assign n1038 = ~g361 & ~g49;
  assign n1039 = ~n1040 & ~n787 & ~n1019;
  assign n1040 = ~g314 & n785;
  assign n1041_1 = g84 & n1042;
  assign n1042 = n1043 & g54 & g59 & g64 & ~n1039 & g79 & g74 & g69;
  assign n1043 = g361 & g49;
  assign n1044 = g84 & ~n1045;
  assign n1045 = ~n1046_1 & ~n1053;
  assign n1046_1 = ~n1047 & n1048 & ~n1052;
  assign n1047 = n1030 & n1048;
  assign n1048 = ~n1049 & ~n1051_1;
  assign n1049 = n778 & n1050;
  assign n1050 = n1019 & ~g301 & ~g310 & ~g319;
  assign n1051_1 = g319 & n778;
  assign n1052 = ~n1037 & ~n1042;
  assign n1053 = ~n1047 & g398 & ~n1048;
  assign n1054 = ~g84 & n1045;
  assign n1055 = ~n785 & ~n1028 & ~n776_1 & ~n787 & ~n1034;
  assign n1056_1 = ~n1057 & ~n1077;
  assign n1057 = n1058 & n1071_1;
  assign n1058 = ~n1059 & ~n1070;
  assign n1059 = n717 & ~n1060;
  assign n1060 = ~n1061_1 & ~n1069;
  assign n1061_1 = n1062 & n1066_1;
  assign n1062 = ~n1063 & ~n1065;
  assign n1063 = g32 & ~n1064;
  assign n1064 = g32 & g36;
  assign n1065 = g36 & ~n1064;
  assign n1066_1 = ~n1067 & ~n1068;
  assign n1067 = g38 & ~g37;
  assign n1068 = ~g38 & g37;
  assign n1069 = ~n1062 & ~n1066_1;
  assign n1070 = ~n717 & n1060;
  assign n1071_1 = ~n1072 & ~n1076_1;
  assign n1072 = g48 & ~n1073;
  assign n1073 = ~n1074 & ~n1075;
  assign n1074 = g39 & ~g40;
  assign n1075 = ~g39 & g40;
  assign n1076_1 = ~g48 & n1073;
  assign n1077 = ~n1058 & ~n1071_1;
  assign n226 = g639 & ~n1079 & ~n1084;
  assign n1079 = g622 & n1080;
  assign n1080 = g619 & n1081_1;
  assign n1081_1 = g616 & n1082;
  assign n1082 = g613 & n1083;
  assign n1083 = g602 & g610;
  assign n1084 = ~g622 & ~n1080;
  assign n231 = g114 | n1086_1;
  assign n1086_1 = n812 & ~n1087;
  assign n1087 = ~g94 & g102;
  assign n1088 = ~n1089 & ~n1095;
  assign n1089 = ~n1094 & ~n1092 & g269 & n1090;
  assign n1090 = ~n931_1 & n1091_1;
  assign n1091_1 = ~n913 & ~n930;
  assign n1092 = g278 & n1093;
  assign n1093 = g276 & g277;
  assign n1094 = ~g278 & ~n1093;
  assign n1095 = ~g269 & g692;
  assign n241 = n1097 | n1098 | ~n1099;
  assign n1097 = g128 & ~g114;
  assign n1098 = ~g128 & g114;
  assign n1099 = ~n806_1 & ~n808;
  assign n246 = g638 & ~n1101_1;
  assign n1101_1 = ~n1102 & ~n1103;
  assign n1102 = g567 & ~n873;
  assign n1103 = g598 & ~n873;
  assign n251 = n1105 | n1106_1;
  assign n1105 = g554 & ~n988;
  assign n1106_1 = ~n911_1 & n988;
  assign n256 = g496 | n1108;
  assign n1108 = ~n1109 & g211 & g210;
  assign n1109 = ~n1110 & ~n1131_1;
  assign n1110 = n970 & ~n1111_1;
  assign n1111_1 = ~n1112 & ~n1130;
  assign n1112 = g471 & ~n1113;
  assign n1113 = ~n1114 & ~n1122;
  assign n1114 = g206 & ~n1115;
  assign n1115 = ~n1116_1 & ~n1119;
  assign n1116_1 = ~g205 & ~n1117 & ~n1118;
  assign n1117 = g693 & ~g204;
  assign n1118 = g204 & g692;
  assign n1119 = g205 & ~n1120 & ~n1121_1;
  assign n1120 = ~g204 & g691;
  assign n1121_1 = g690 & g204;
  assign n1122 = ~g206 & ~n1123;
  assign n1123 = ~n1124 & ~n1127;
  assign n1124 = ~g205 & ~n1125 & ~n1126_1;
  assign n1125 = g697 & ~g204;
  assign n1126_1 = g696 & g204;
  assign n1127 = g205 & ~n1128 & ~n1129;
  assign n1128 = g695 & ~g204;
  assign n1129 = g204 & g694;
  assign n1130 = ~g471 & n1113;
  assign n1131_1 = ~n970 & ~n1132;
  assign n1132 = ~n978 & ~n1133;
  assign n1133 = g471 & ~n1134;
  assign n1134 = g471 & n967;
  assign n261 = n1136_1 | n1166_1;
  assign n1136_1 = n1137 & ~n1155 & ~n1165;
  assign n1137 = ~n806_1 & ~n1138;
  assign n1138 = ~n1139 & ~n1144;
  assign n1139 = ~n1140 & ~n1142;
  assign n1140 = n807 & ~n1141_1;
  assign n1141_1 = ~g94 & ~g98;
  assign n1142 = n808 & n1143;
  assign n1143 = ~g107 & g89 & g102;
  assign n1144 = ~n1145 & ~n1151_1;
  assign n1145 = ~g188 & n1146_1;
  assign n1146_1 = ~g179 & n1147;
  assign n1147 = n1149 & ~g170 & ~g161 & n1148;
  assign n1148 = ~g143 & ~g152;
  assign n1149 = ~n1150 & ~n816_1 & ~n1087;
  assign n1150 = ~g102 & n814;
  assign n1151_1 = g188 & n1152;
  assign n1152 = g179 & n1153;
  assign n1153 = ~n1149 & g170 & g161 & n1154;
  assign n1154 = g143 & g152;
  assign n1155 = g179 & ~n1156_1;
  assign n1156_1 = ~n1157 & ~n1164;
  assign n1157 = ~n1158 & n1159 & ~n1163;
  assign n1158 = n1139 & n1159;
  assign n1159 = ~n1160 & ~n1162;
  assign n1160 = n808 & n1161_1;
  assign n1161_1 = n1087 & ~g89 & ~g98 & ~g107;
  assign n1162 = g107 & n808;
  assign n1163 = ~n1147 & ~n1153;
  assign n1164 = ~n1158 & g184 & ~n1159;
  assign n1165 = ~g179 & n1156_1;
  assign n1166_1 = ~n814 & ~n1137 & ~n806_1 & ~n816_1 & ~n1143;
  assign n271 = ~n1168 | n1178;
  assign n1168 = g639 & ~n1169;
  assign n1169 = g594 & n1170;
  assign n1170 = g590 & n1171_1;
  assign n1171_1 = g574 & n1172;
  assign n1172 = g586 & n1173;
  assign n1173 = g582 & n1174;
  assign n1174 = g578 & n1175;
  assign n1175 = g631 & n1176_1;
  assign n1176_1 = g628 & n1177;
  assign n1177 = g625 & n1079;
  assign n1178 = ~n1170 & ~n1179;
  assign n1179 = ~g590 & ~n1171_1;
  assign n276 = n1181_1 | n1182;
  assign n1181_1 = g551 & ~n988;
  assign n1182 = ~n961_1 & n988;
  assign n286 = n1206 | n1203 | n1184 | n1190 | n1202 | n1204 | n1208 | n1209 | n1211 | n1215 | n1222 | n1224 | n1226;
  assign n1184 = g562 & n1185;
  assign n1185 = n1187 & g678 & n1186_1 & ~g680 & g679;
  assign n1186_1 = g698 & g688 & g689;
  assign n1187 = ~n1188 & g699 & g41 & g702;
  assign n1188 = ~n794 & ~n1189;
  assign n1189 = ~g658 & g266;
  assign n1190 = ~n1201_1 & ~n1200 & ~n1199 & ~n1198 & ~n1197 & ~n1194 & ~n801_1 & ~n1185 & ~n1191_1 & ~n1192 & ~n1193 & n1196_1;
  assign n1191_1 = n1187 & n1024 & ~g683 & g684;
  assign n1192 = n793 & n821_1 & ~g684 & ~g685;
  assign n1193 = ~g688 & n793 & n861_1;
  assign n1194 = n1195 & n1024 & g682;
  assign n1195 = n1187 & g684 & g683;
  assign n1196_1 = ~n792 & ~n820;
  assign n1197 = ~g679 & n1187 & n1186_1 & g678 & ~g680;
  assign n1198 = n1195 & n1024 & ~g682 & ~g681;
  assign n1199 = ~g680 & ~g679 & n1186_1 & ~g678 & n1187;
  assign n1200 = n1187 & g680 & n1186_1 & ~g678 & ~g679;
  assign n1201_1 = g681 & ~g682 & n1195 & n1024;
  assign n1202 = g293 & n1191_1;
  assign n1203 = g551 & n1201_1;
  assign n1204 = g508 & n1205;
  assign n1205 = g677 & n1198;
  assign n1206 = g536 & n1207;
  assign n1207 = ~g677 & n1198;
  assign n1208 = g692 & n1192;
  assign n1209 = ~n1088 & n1210;
  assign n1210 = g687 & n1193;
  assign n1211 = n801_1 & ~n1212;
  assign n1212 = ~n1213 & ~n1214;
  assign n1213 = ~g677 & g692;
  assign n1214 = g677 & g692;
  assign n1215 = ~n1216 & n1221;
  assign n1216 = ~n1217 & ~n1220;
  assign n1217 = ~n1219 & ~n981_1 & g197 & n1218;
  assign n1218 = ~n966_1 & n975;
  assign n1219 = ~g206 & ~n982;
  assign n1220 = ~g197 & g692;
  assign n1221 = ~g687 & n1193;
  assign n1222 = g453 & n1223;
  assign n1223 = ~g677 & n1194;
  assign n1224 = g410 & n1225;
  assign n1225 = g677 & n1194;
  assign n1226 = g692 & ~n1196_1;
  assign n291 = g638 & ~n1228 & ~n1230;
  assign n1228 = g606 & n1229;
  assign n1229 = g642 & n881_1;
  assign n1230 = ~g606 & ~n1229;
  assign n296 = n1166_1 | n1232;
  assign n1232 = n1137 & ~n1233 & ~n1238;
  assign n1233 = g188 & ~n1234;
  assign n1234 = ~n1235 & ~n1237;
  assign n1235 = ~n1158 & n1159 & ~n1236;
  assign n1236 = ~n1146_1 & ~n1152;
  assign n1237 = ~n1158 & g193 & ~n1159;
  assign n1238 = ~g188 & n1234;
  assign n301 = g638 & ~n1240 & ~n1241;
  assign n1240 = g646 & n1228;
  assign n1241 = ~g646 & ~n1228;
  assign n306 = g326 & ~n1018;
  assign n311 = n1055 | n1244;
  assign n1244 = n1028 & ~n1245 & ~n1249;
  assign n1245 = g361 & ~n1246;
  assign n1246 = ~n1247 & ~n1248;
  assign n1247 = g366 & ~n1047;
  assign n1248 = n1048 & ~n1047;
  assign n1249 = ~g361 & n1246;
  assign n321 = n1251 | n1253;
  assign n1251 = g398 & ~n776_1 & ~n1252;
  assign n1252 = ~g301 & n1051_1;
  assign n1253 = g394 & n1252;
  assign n331 = g639 & ~n1080 & ~n1255;
  assign n1255 = ~g619 & ~n1081_1;
  assign n1256 = ~n1257 & ~n1262;
  assign n1257 = g197 & ~n1258;
  assign n1258 = n1218 & ~n1259;
  assign n1259 = ~n1260 & ~n1261;
  assign n1260 = g208 & n980;
  assign n1261 = ~g208 & ~n980;
  assign n1262 = ~g197 & g694;
  assign n346 = n1264 | n1265;
  assign n1264 = ~n1252 & g390 & ~n776_1;
  assign n1265 = g386 & n1252;
  assign n351 = g639 & ~n1177 & ~n1267;
  assign n1267 = ~g625 & ~n1079;
  assign n361 = n1269 | n1270;
  assign n1269 = g437 & ~n987;
  assign n1270 = g441 & n987;
  assign n1271 = ~n1272 & ~n1273;
  assign n1272 = g269 & ~g276 & n1090;
  assign n1273 = ~g269 & g690;
  assign n371 = n1279 | n1277 | n1190 | n1275 | n1276 | n1278 | n1280 | n1281 | n1282 | n1283 | n1284 | n1285 | n1289 | n1293 | n1294 | n1295;
  assign n1275 = g669 & n1200;
  assign n1276 = g564 & n1185;
  assign n1277 = g545 & n1201_1;
  assign n1278 = g197 & n1191_1;
  assign n1279 = g532 & n1207;
  assign n1280 = g500 & n1205;
  assign n1281 = ~g486 & n1197;
  assign n1282 = g496 & n1199;
  assign n1283 = g690 & n1192;
  assign n1284 = n1210 & ~n1271;
  assign n1285 = n801_1 & ~n1286;
  assign n1286 = ~n1287 & ~n1288;
  assign n1287 = g690 & ~g677;
  assign n1288 = g690 & g677;
  assign n1289 = n1221 & ~n1290;
  assign n1290 = ~n1291 & ~n1292;
  assign n1291 = g197 & ~g204 & n1218;
  assign n1292 = g690 & ~g197;
  assign n1293 = g461 & n1223;
  assign n1294 = g402 & n1225;
  assign n1295 = g690 & ~n1196_1;
  assign n376 = g331 & ~n1018;
  assign n391 = ~n1298 & ~n1300;
  assign n1298 = g582 & g586 & g578 & g574 & n1299;
  assign n1299 = ~g590 & g594;
  assign n1300 = ~n1315 & ~n1301 & ~n1308 & ~n1299;
  assign n1301 = ~g586 & ~n1302 & ~n1305;
  assign n1302 = ~g582 & ~n1303 & ~n1304;
  assign n1303 = g697 & ~g578;
  assign n1304 = g696 & g578;
  assign n1305 = g582 & ~n1306 & ~n1307;
  assign n1306 = g695 & ~g578;
  assign n1307 = g578 & g694;
  assign n1308 = g586 & ~n1309 & ~n1312;
  assign n1309 = ~g582 & ~n1310 & ~n1311;
  assign n1310 = g693 & ~g578;
  assign n1311 = g578 & g692;
  assign n1312 = g582 & ~n1313 & ~n1314;
  assign n1313 = ~g578 & g691;
  assign n1314 = g690 & g578;
  assign n1315 = g590 & ~g594;
  assign n396 = n1317 | n1319;
  assign n1317 = g157 & ~n806_1 & ~n1318;
  assign n1318 = ~g89 & n1162;
  assign n1319 = g148 & n1318;
  assign n1320 = ~n1321 & ~n1322;
  assign n1321 = g269 & ~n961_1;
  assign n1322 = ~g269 & g696;
  assign n416 = n1324 | n1325;
  assign n1324 = g449 & ~n987;
  assign n1325 = g453 & n987;
  assign n421 = g117 & ~n1086_1;
  assign n426 = n1328 | n1330;
  assign n1328 = g528 & ~n1329;
  assign n1329 = g677 & n1023;
  assign n1330 = g697 & n1329;
  assign n436 = n1332 | n1333;
  assign n1332 = g426 & ~n987;
  assign n1333 = g422 & n987;
  assign n441 = g638 & ~n881_1 & ~n1335;
  assign n1335 = ~g634 & ~n873;
  assign n446 = g669 | n1337;
  assign n1337 = ~g22 & n1056_1;
  assign n451 = n1339 | n1340;
  assign n1339 = g520 & ~n1329;
  assign n1340 = g695 & n1329;
  assign n1341 = ~n1342 & ~n1348;
  assign n1342 = ~n1343 & g269 & n1091_1;
  assign n1343 = ~n931_1 & ~n1344 & ~n1347;
  assign n1344 = g281 & ~n1345;
  assign n1345 = g280 & n1346;
  assign n1346 = g279 & n1092;
  assign n1347 = ~g281 & n1345;
  assign n1348 = g695 & ~g269;
  assign n461 = n1350 | n1351;
  assign n1350 = ~n1318 & g175 & ~n806_1;
  assign n1351 = g166 & n1318;
  assign n466 = n1357 | n1355 | n1190 | n1353 | n1354 | n1356 | n1358 | n1359 | n1366 | n1370 | n1371 | n1372 | n1373;
  assign n1353 = g561 & n1185;
  assign n1354 = g297 & n1191_1;
  assign n1355 = g554 & n1201_1;
  assign n1356 = g512 & n1205;
  assign n1357 = g541 & n1207;
  assign n1358 = g693 & n1192;
  assign n1359 = n1210 & ~n1360;
  assign n1360 = ~n1361 & ~n1365;
  assign n1361 = g269 & ~n931_1 & ~n1362;
  assign n1362 = n1091_1 & ~n1363;
  assign n1363 = ~n1346 & ~n1364;
  assign n1364 = ~g279 & ~n1092;
  assign n1365 = g693 & ~g269;
  assign n1366 = n801_1 & ~n1367;
  assign n1367 = ~n1368 & ~n1369;
  assign n1368 = g693 & ~g677;
  assign n1369 = g693 & g677;
  assign n1370 = ~n964 & n1221;
  assign n1371 = g449 & n1223;
  assign n1372 = g414 & n1225;
  assign n1373 = g693 & ~n1196_1;
  assign n471 = g639 & ~n1175 & ~n1375;
  assign n1375 = ~g631 & ~n1176_1;
  assign n476 = n1055 | n1377;
  assign n1377 = n1028 & ~n1378 & ~n1385;
  assign n1378 = g69 & ~n1379;
  assign n1379 = ~n1380 & ~n1384;
  assign n1380 = ~n1047 & n1048 & ~n1381;
  assign n1381 = ~n1382 & ~n1383;
  assign n1382 = n1039 & n1038 & ~g64 & ~g59 & ~g54;
  assign n1383 = n1043 & ~n1039 & g64 & g59 & g54;
  assign n1384 = ~n1047 & g386 & ~n1048;
  assign n1385 = ~g69 & n1379;
  assign n486 = g301 & ~g314;
  assign n491 = n1388 | n1389;
  assign n1388 = g457 & ~n987;
  assign n1389 = g461 & n987;
  assign n506 = g327 & ~n1018;
  assign n516 = n1392 | n1393;
  assign n1392 = g418 & ~n987;
  assign n1393 = g414 & n987;
  assign n521 = n1395 | n1396;
  assign n1395 = g402 & ~n987;
  assign n1396 = n987 & ~n1397;
  assign n1397 = ~n1398 & ~n1399;
  assign n1398 = ~g465 & g471;
  assign n1399 = g465 & g478;
  assign n526 = n1401 | n1403;
  assign n1401 = g297 & ~n1402;
  assign n1402 = n799 & n1024 & ~g683 & g684;
  assign n1403 = g693 & n1402;
  assign n536 = n1405 | n1406;
  assign n1405 = g410 & ~n987;
  assign n1406 = g406 & n987;
  assign n541 = n1408 | n1409;
  assign n1408 = g430 & ~n987;
  assign n1409 = g426 & n987;
  assign n546 = n1418 | n1413 | n1190 | n1411 | n1412 | n1414 | n1422 | n1437 | n1438 | n1439;
  assign n1411 = g528 & n1205;
  assign n1412 = g557 & n1185;
  assign n1413 = g697 & n1192;
  assign n1414 = n1210 & ~n1415;
  assign n1415 = ~n1416 & ~n1417;
  assign n1416 = g269 & ~n911_1;
  assign n1417 = g697 & ~g269;
  assign n1418 = n801_1 & ~n1419;
  assign n1419 = ~n1420 & ~n1421;
  assign n1420 = g697 & ~g677;
  assign n1421 = g697 & g677;
  assign n1422 = n1221 & ~n1423;
  assign n1423 = ~n1424 & ~n1436;
  assign n1424 = g197 & ~n1425;
  assign n1425 = ~n1426 & ~n1434 & ~n1435;
  assign n1426 = ~n1429 & ~n966_1 & ~n977 & ~n1427 & g211;
  assign n1427 = n1131_1 & n1428;
  assign n1428 = ~g211 & g210;
  assign n1429 = n976_1 & ~n1430;
  assign n1430 = ~n1431 & n1432;
  assign n1431 = g211 & ~g210;
  assign n1432 = ~n1108 & ~n1433;
  assign n1433 = n1110 & n1428;
  assign n1434 = ~n1433 & n976_1 & n1428;
  assign n1435 = ~n976_1 & ~n1432;
  assign n1436 = g697 & ~g197;
  assign n1437 = g434 & n1223;
  assign n1438 = g430 & n1225;
  assign n1439 = g697 & ~n1196_1;
  assign n556 = n1441 | n1442;
  assign n1441 = g453 & ~n987;
  assign n1442 = g457 & n987;
  assign n561 = n1444 | n1445;
  assign n1444 = g269 & ~n1402;
  assign n1445 = g691 & n1402;
  assign n566 = ~n1168 | n1447;
  assign n1447 = ~n1171_1 & ~n1448;
  assign n1448 = ~g574 & ~n1172;
  assign n571 = n1450 | n1451;
  assign n1450 = g441 & ~n987;
  assign n1451 = g445 & n987;
  assign n581 = ~n1453 | n1454 | n1456;
  assign n1453 = ~n776_1 & ~n778;
  assign n1454 = g349 & ~n1455;
  assign n1455 = g323 & n780;
  assign n1456 = ~g349 & n1455;
  assign n591 = n1168 & ~n1172 & ~n1458;
  assign n1458 = ~g586 & ~n1173;
  assign n596 = g638 & ~n1460 & ~n1463;
  assign n1460 = g571 & n1461;
  assign n1461 = g654 & n1462;
  assign n1462 = g650 & n1240;
  assign n1463 = ~g571 & ~n1461;
  assign n601 = n1469 | n1467 | n1190 | n1465 | n1466 | n1468 | n1473 | n1479 | n1480 | n1481;
  assign n1465 = g524 & n1205;
  assign n1466 = g558 & n1185;
  assign n1467 = g696 & n1192;
  assign n1468 = n1210 & ~n1320;
  assign n1469 = n801_1 & ~n1470;
  assign n1470 = ~n1471 & ~n1472;
  assign n1471 = g696 & ~g677;
  assign n1472 = g696 & g677;
  assign n1473 = n1221 & ~n1474;
  assign n1474 = ~n1475 & ~n1478;
  assign n1475 = g197 & ~n1476;
  assign n1476 = ~n1434 & ~n1477 & ~n966_1 & ~n1429;
  assign n1477 = ~n1435 & ~n977 & ~n1427 & g210;
  assign n1478 = g696 & ~g197;
  assign n1479 = g437 & n1223;
  assign n1480 = g426 & n1225;
  assign n1481 = g696 & ~n1196_1;
  assign n606 = g323 | n1018;
  assign n616 = g638 & ~n1461 & ~n1484;
  assign n1484 = ~g654 & ~n1462;
  assign n621 = n1486 | n1487;
  assign n1486 = g293 & ~n1402;
  assign n1487 = g692 & n1402;
  assign n631 = n1489 | n1490;
  assign n1489 = g445 & ~n987;
  assign n1490 = g449 & n987;
  assign n636 = n1492 | n1493;
  assign n1492 = ~n1252 & g374 & ~n776_1;
  assign n1493 = g370 & n1252;
  assign n651 = ~n1453 | n1495;
  assign n1495 = g357 & ~n1496;
  assign n1496 = g323 & n779;
  assign n656 = n1498 | n1499;
  assign n1498 = ~n1252 & g386 & ~n776_1;
  assign n1499 = g382 & n1252;
  assign n661 = n1501 | n1502;
  assign n1501 = g504 & ~n1329;
  assign n1502 = g691 & n1329;
  assign n671 = n1504 | n1505;
  assign n1504 = ~n1318 & g166 & ~n806_1;
  assign n1505 = g157 & n1318;
  assign n676 = n1507 | n1513;
  assign n1507 = ~n1022 & ~n1508;
  assign n1508 = ~g541 & ~n1509;
  assign n1509 = ~g536 & n988 & ~n1510;
  assign n1510 = ~n1511 & ~n1512;
  assign n1511 = ~g465 & n976_1;
  assign n1512 = g465 & n930;
  assign n1513 = g693 & n1022;
  assign n681 = n1055 | n1515;
  assign n1515 = n1028 & ~n1516 & ~n1523;
  assign n1516 = g74 & ~n1517;
  assign n1517 = ~n1518 & ~n1522;
  assign n1518 = ~n1047 & n1048 & ~n1519;
  assign n1519 = ~n1520 & ~n1521;
  assign n1520 = n1039 & ~g54 & ~g69 & ~g64 & ~g59 & n1038;
  assign n1521 = n1043 & g54 & ~n1039 & g69 & g64 & g59;
  assign n1522 = ~n1047 & g390 & ~n1048;
  assign n1523 = ~g74 & n1517;
  assign n686 = ~n1453 | n1525 | n1526;
  assign n1525 = ~g323 & g338;
  assign n1526 = g323 & ~g338;
  assign n696 = n1528 | n1529;
  assign n1528 = g516 & ~n1329;
  assign n1529 = g694 & n1329;
  assign n701 = n1531 | n1535;
  assign n1531 = ~n1022 & g536 & ~n1532;
  assign n1532 = n988 & ~n1533 & ~n1534;
  assign n1533 = ~g465 & ~n968;
  assign n1534 = g465 & ~n920;
  assign n1535 = g692 & n1022;
  assign n711 = n1453 & ~n1537 & ~n1538;
  assign n1537 = ~g353 & ~n1456;
  assign n1538 = g353 & n1456;
  assign n716 = n1540 | n1541;
  assign n1540 = g545 & ~n988;
  assign n1541 = n988 & ~n1476;
  assign n726 = ~n1453 | n1543 | n1544;
  assign n1543 = g341 & ~n1526;
  assign n1544 = ~g341 & n1526;
  assign n746 = n1546 | n1557;
  assign n1546 = ~n776_1 & ~n1547;
  assign n1547 = ~n787 & ~n1548;
  assign n1548 = g336 & ~n1549;
  assign n1549 = ~n1556 & ~n1552 & ~n486 & g328 & ~n1550;
  assign n1550 = ~n1050 & ~n1551 & ~n785 & ~n1034 & ~n784 & ~n786_1;
  assign n1551 = g301 & g319;
  assign n1552 = n1415 & ~n1553;
  assign n1553 = ~n1554 & ~n1555;
  assign n1554 = g332 & ~n786_1;
  assign n1555 = ~n1034 & ~g332 & ~n1551 & ~n784;
  assign n1556 = ~n1415 & n1553;
  assign n1557 = n776_1 & ~n1558;
  assign n1558 = ~n1559 & ~n1585 & ~n1646;
  assign n1559 = ~n1560 & ~n1572;
  assign n1560 = ~n1561 & ~n1566;
  assign n1561 = ~n1562 & ~n1565;
  assign n1562 = g269 & ~n1563;
  assign n1563 = ~n836_1 & ~n1564;
  assign n1564 = g230 & ~g658;
  assign n1565 = g681 & ~g269;
  assign n1566 = ~n1567 & ~n1571;
  assign n1567 = g269 & ~n1568;
  assign n1568 = ~n1569 & ~n1570;
  assign n1569 = g634 & g658;
  assign n1570 = g224 & ~g658;
  assign n1571 = ~g269 & g680;
  assign n1572 = ~n1573 & ~n1579;
  assign n1573 = ~n1574 & ~n1578;
  assign n1574 = g269 & ~n1575;
  assign n1575 = ~n1576 & ~n1577;
  assign n1576 = g598 & g658;
  assign n1577 = g218 & ~g658;
  assign n1578 = ~g269 & g679;
  assign n1579 = ~n1580 & ~n1584;
  assign n1580 = g269 & ~n1581;
  assign n1581 = ~n1582 & ~n1583;
  assign n1582 = g567 & g658;
  assign n1583 = g212 & ~g658;
  assign n1584 = g678 & ~g269;
  assign n1585 = ~n1586 & ~n1591;
  assign n1586 = ~g337 & ~n1587;
  assign n1587 = ~n1590 & ~n1210 & ~n1588 & ~n1589;
  assign n1588 = g269 & n791_1;
  assign n1589 = g269 & n794;
  assign n1590 = n803 & ~g269 & n861_1 & ~g688;
  assign n1591 = ~n1592 & ~n1643;
  assign n1592 = ~n1593 & ~n1608 & ~n1619;
  assign n1593 = ~n1594 & ~n1601;
  assign n1594 = ~n1595 & ~n1598;
  assign n1595 = ~n1596 & ~n1597;
  assign n1596 = g197 & ~n1563;
  assign n1597 = g681 & ~g197;
  assign n1598 = ~n1599 & ~n1600;
  assign n1599 = g197 & ~n1568;
  assign n1600 = g680 & ~g197;
  assign n1601 = ~n1602 & ~n1605;
  assign n1602 = ~n1603 & ~n1604;
  assign n1603 = g197 & ~n1575;
  assign n1604 = g679 & ~g197;
  assign n1605 = ~n1606 & ~n1607;
  assign n1606 = g197 & ~n1581;
  assign n1607 = g678 & ~g197;
  assign n1608 = ~n1609 & ~n1614 & ~n1618;
  assign n1609 = ~g337 & ~n1610;
  assign n1610 = ~n1613 & ~n1221 & ~n1611 & ~n1612;
  assign n1611 = g197 & n791_1;
  assign n1612 = g197 & n794;
  assign n1613 = n797 & ~g197 & n861_1 & ~g688;
  assign n1614 = g197 & ~n1615;
  assign n1615 = ~n1616 & ~n1617;
  assign n1616 = g571 & g658;
  assign n1617 = ~g658 & g260;
  assign n1618 = g686 & ~g197;
  assign n1619 = ~n1620 & ~n1632;
  assign n1620 = ~n1621 & ~n1627;
  assign n1621 = ~n1622 & ~n1626;
  assign n1622 = g197 & ~n1623;
  assign n1623 = ~n1624 & ~n1625;
  assign n1624 = g654 & g658;
  assign n1625 = g254 & ~g658;
  assign n1626 = g685 & ~g197;
  assign n1627 = ~n1628 & ~n1631;
  assign n1628 = g197 & ~n1629;
  assign n1629 = ~n826_1 & ~n1630;
  assign n1630 = g248 & ~g658;
  assign n1631 = g684 & ~g197;
  assign n1632 = ~n1633 & ~n1638;
  assign n1633 = ~n1634 & ~n1637;
  assign n1634 = g197 & ~n1635;
  assign n1635 = ~n829 & ~n1636;
  assign n1636 = g242 & ~g658;
  assign n1637 = g683 & ~g197;
  assign n1638 = ~n1639 & ~n1642;
  assign n1639 = g197 & ~n1640;
  assign n1640 = ~n833 & ~n1641;
  assign n1641 = ~g658 & g236;
  assign n1642 = g682 & ~g197;
  assign n1643 = ~n1644 & ~n1645;
  assign n1644 = g269 & ~n1615;
  assign n1645 = ~g269 & g686;
  assign n1646 = ~n1647 & ~n1654;
  assign n1647 = ~n1648 & ~n1651;
  assign n1648 = ~n1649 & ~n1650;
  assign n1649 = g269 & ~n1623;
  assign n1650 = g685 & ~g269;
  assign n1651 = ~n1652 & ~n1653;
  assign n1652 = g269 & ~n1629;
  assign n1653 = g684 & ~g269;
  assign n1654 = ~n1655 & ~n1658;
  assign n1655 = ~n1656 & ~n1657;
  assign n1656 = g269 & ~n1635;
  assign n1657 = ~g269 & g683;
  assign n1658 = ~n1659 & ~n1660;
  assign n1659 = g269 & ~n1640;
  assign n1660 = g682 & ~g269;
  assign n751 = ~n1453 | n1662 | n1663;
  assign n1662 = g345 & ~n1544;
  assign n1663 = ~g345 & n1544;
  assign n756 = g639 & ~n1176_1 & ~n1665;
  assign n1665 = ~g628 & ~n1177;
  assign n781 = ~g639 | n1667;
  assign n1667 = g639 & ~n1082 & ~n1668;
  assign n1668 = ~g613 & ~n1083;
  assign n801 = n1166_1 | n1670;
  assign n1670 = n1137 & ~n1671 & ~n1675;
  assign n1671 = g143 & ~n1672;
  assign n1672 = ~n1673 & ~n1674;
  assign n1673 = g148 & ~n1158;
  assign n1674 = n1159 & ~n1158;
  assign n1675 = ~g143 & n1672;
  assign n806 = g672 | n1677;
  assign n1677 = ~g22 & n714;
  assign n816 = n1679 | n776_1 | n1680;
  assign n1679 = g398 & n1252;
  assign n1680 = g366 & ~n1252;
  assign n826 = g492 | n956_1;
  assign n831 = n1166_1 | n1683;
  assign n1683 = n1137 & ~n1684 & ~n1691;
  assign n1684 = g170 & ~n1685;
  assign n1685 = ~n1686 & ~n1690;
  assign n1686 = ~n1158 & n1159 & ~n1687;
  assign n1687 = ~n1688 & ~n1689;
  assign n1688 = ~g161 & n1148 & n1149;
  assign n1689 = ~n1149 & g161 & n1154;
  assign n1690 = ~n1158 & g175 & ~n1159;
  assign n1691 = ~g170 & n1685;
  assign n851 = g639 & ~g602;
  assign n856 = g638 & ~n1229 & ~n1694;
  assign n1694 = ~g642 & ~n881_1;
  assign n1695 = ~n1696 & ~n1700;
  assign n1696 = g269 & ~n1697;
  assign n1697 = n1090 & ~n1698;
  assign n1698 = ~n1345 & ~n1699;
  assign n1699 = ~g280 & ~n1346;
  assign n1700 = ~g269 & g694;
  assign n871 = g639 & ~n1702;
  assign n1702 = ~n1703 & ~n1704;
  assign n1703 = g602 & ~n1083;
  assign n1704 = g610 & ~n1083;
  assign n876 = n1706 | n806_1 | n1707;
  assign n1706 = g193 & n1318;
  assign n1707 = g148 & ~n1318;
  assign n1708 = ~n1709 & ~n1713;
  assign n1709 = ~n1710 & g197 & n975;
  assign n1710 = ~n966_1 & ~n1711 & ~n1712;
  assign n1711 = g209 & ~n1260;
  assign n1712 = ~g209 & n1260;
  assign n1713 = g695 & ~g197;
  assign n896 = g119 & ~n1086_1;
  assign n901 = n1055 | n1716;
  assign n1716 = n1028 & ~n1717 & ~n1725;
  assign n1717 = g54 & ~n1718;
  assign n1718 = ~n1719 & ~n1720;
  assign n1719 = ~n1047 & g374 & ~n1048;
  assign n1720 = ~n1724 & ~n1047 & n1048 & ~n1721;
  assign n1721 = ~n1722 & ~n1723;
  assign n1722 = ~g361 & n1039;
  assign n1723 = g361 & ~n1039;
  assign n1724 = ~n1038 & ~n1043;
  assign n1725 = ~g54 & n1718;
  assign n906 = n1168 & ~n1169 & ~n1727;
  assign n1727 = ~g594 & ~n1170;
  assign n921 = g639 & ~n1081_1 & ~n1729;
  assign n1729 = ~g616 & ~n1082;
  assign n926 = n1055 | n1731;
  assign n1731 = n1028 & ~n1732 & ~n1739;
  assign n1732 = g79 & ~n1733;
  assign n1733 = ~n1734 & ~n1738;
  assign n1734 = ~n1047 & n1048 & ~n1735;
  assign n1735 = ~n1736 & ~n1737;
  assign n1736 = n1039 & n1038 & ~g59 & ~g74 & ~g69 & ~g64 & ~g54;
  assign n1737 = n1043 & g54 & g59 & ~n1039 & g74 & g69 & g64;
  assign n1738 = ~n1047 & g394 & ~n1048;
  assign n1739 = ~g79 & n1733;
  assign n941 = n1168 & ~n1174 & ~n1741;
  assign n1741 = ~g578 & ~n1175;
  assign n946 = n1743 | n1744;
  assign n1743 = ~n1318 & g184 & ~n806_1;
  assign n1744 = g175 & n1318;
  assign n951 = g118 & ~n1086_1;
  assign n1746 = ~n1425 & ~n1476;
  assign n961 = ~n1099 | n1748;
  assign n1748 = g139 & ~n1749;
  assign n1749 = g114 & n809;
  assign n966 = n1751 | n1752;
  assign n1751 = g422 & ~n987;
  assign n1752 = g418 & n987;
  assign n976 = n1754 | n1755;
  assign n1754 = ~n1252 & g394 & ~n776_1;
  assign n1755 = g390 & n1252;
  assign n986 = n1761 | n1759 | n1190 | n1757 | n1758 | n1760 | n1765 | n1766 | n1767 | n1768;
  assign n1757 = g520 & n1205;
  assign n1758 = g559 & n1185;
  assign n1759 = g695 & n1192;
  assign n1760 = n1210 & ~n1341;
  assign n1761 = n801_1 & ~n1762;
  assign n1762 = ~n1763 & ~n1764;
  assign n1763 = g695 & ~g677;
  assign n1764 = g695 & g677;
  assign n1765 = n1221 & ~n1708;
  assign n1766 = g441 & n1223;
  assign n1767 = g422 & n1225;
  assign n1768 = g695 & ~n1196_1;
  assign n996 = g45 & ~g658;
  assign n1001 = g638 & ~n1462 & ~n1771;
  assign n1771 = ~g650 & ~n1240;
  assign n1006 = n1773 | n1774;
  assign n1773 = ~n1252 & g378 & ~n776_1;
  assign n1774 = g374 & n1252;
  assign n1011 = n1776 | n1777;
  assign n1776 = g508 & ~n1329;
  assign n1777 = g692 & n1329;
  assign n1016 = n1779 | n1780;
  assign n1779 = g548 & ~n988;
  assign n1780 = n988 & ~n1425;
  assign n1021 = n1782 | n1783;
  assign n1782 = ~n1252 & g370 & ~n776_1;
  assign n1783 = g366 & n1252;
  assign n1026 = n1785 | n1786;
  assign n1785 = g406 & ~n987;
  assign n1786 = g402 & n987;
  assign n1036 = n1788 | n1789;
  assign n1788 = g500 & ~n1329;
  assign n1789 = g690 & n1329;
  assign n1790 = ~n1791 & ~n1795;
  assign n1791 = ~n1792 & g197 & n1218;
  assign n1792 = ~n1793 & ~n1794;
  assign n1793 = g204 & ~n982;
  assign n1794 = g205 & ~n982;
  assign n1795 = ~g197 & g691;
  assign n1046 = n1797 | n1798;
  assign n1797 = g197 & ~n1402;
  assign n1798 = g690 & n1402;
  assign n1056 = g122 & ~n1086_1;
  assign n1061 = n1801 | n1802;
  assign n1801 = g524 & ~n1329;
  assign n1802 = g696 & n1329;
  assign n1071 = ~n806_1 & ~n1804 & ~n1806;
  assign n1804 = g111 & n1805;
  assign n1805 = n1143 & n1138;
  assign n1806 = ~g111 & ~n1805;
  assign n1076 = ~n1099 | n1808 | n1809;
  assign n1808 = g131 & ~n1098;
  assign n1809 = ~g131 & n1098;
  assign n1081 = n1815 | n1813 | n1190 | n1811 | n1812 | n1814 | n1816 | n1817 | n1818 | n1819 | n1820 | n1827 | n1831 | n1832 | n1833 | n1834;
  assign n1811 = g672 & n1200;
  assign n1812 = g563 & n1185;
  assign n1813 = g548 & n1201_1;
  assign n1814 = g269 & n1191_1;
  assign n1815 = g465 & n1207;
  assign n1816 = g504 & n1205;
  assign n1817 = ~g489 & n1197;
  assign n1818 = g492 & n1199;
  assign n1819 = g691 & n1192;
  assign n1820 = n1210 & ~n1821;
  assign n1821 = ~n1822 & ~n1826;
  assign n1822 = ~n1823 & g269 & n1090;
  assign n1823 = ~n1824 & ~n1825;
  assign n1824 = g276 & ~n1093;
  assign n1825 = g277 & ~n1093;
  assign n1826 = ~g269 & g691;
  assign n1827 = n801_1 & ~n1828;
  assign n1828 = ~n1829 & ~n1830;
  assign n1829 = ~g677 & g691;
  assign n1830 = g677 & g691;
  assign n1831 = n1221 & ~n1790;
  assign n1832 = g457 & n1223;
  assign n1833 = g406 & n1225;
  assign n1834 = g691 & ~n1196_1;
  assign n1086 = n1840 | n1838 | n1190 | n1836 | n1837 | n1839 | n1844 | n1845 | n1846 | n1847;
  assign n1836 = g516 & n1205;
  assign n1837 = g560 & n1185;
  assign n1838 = g694 & n1192;
  assign n1839 = n1210 & ~n1695;
  assign n1840 = n801_1 & ~n1841;
  assign n1841 = ~n1842 & ~n1843;
  assign n1842 = ~g677 & g694;
  assign n1843 = g677 & g694;
  assign n1844 = n1221 & ~n1256;
  assign n1845 = g445 & n1223;
  assign n1846 = g418 & n1225;
  assign n1847 = g694 & ~n1196_1;
  assign n1096 = n1168 & ~n1173 & ~n1849;
  assign n1849 = ~g582 & ~n1174;
  assign n1111 = n1851 | n1852;
  assign n1851 = ~n1318 & g193 & ~n806_1;
  assign n1852 = g184 & n1318;
  assign n1116 = ~n1099 | n1854 | n1855;
  assign n1854 = g135 & ~n1809;
  assign n1855 = ~g135 & n1809;
  assign n1121 = n1857 | n1858;
  assign n1857 = ~n1252 & g382 & ~n776_1;
  assign n1858 = g378 & n1252;
  assign n1126 = n1860 | n1861;
  assign n1860 = g414 & ~n987;
  assign n1861 = g410 & n987;
  assign n1131 = n1863 | n1864;
  assign n1863 = g434 & ~n987;
  assign n1864 = g437 & n987;
  assign n1136 = g45 & ~g266;
  assign n1141 = n1055 | n1867;
  assign n1867 = n1028 & ~n1868 & ~n1872;
  assign n1868 = g49 & ~n1869;
  assign n1869 = ~n1870 & ~n1871;
  assign n1870 = ~n1047 & n1048 & ~n1721;
  assign n1871 = ~n1047 & g370 & ~n1048;
  assign n1872 = ~g49 & n1869;
  assign n1146 = n1166_1 | n1874;
  assign n1874 = n1137 & ~n1875 & ~n1882;
  assign n1875 = g152 & ~n1876;
  assign n1876 = ~n1877 & ~n1881;
  assign n1877 = ~n1158 & n1159 & ~n1878;
  assign n1878 = ~n1879 & ~n1880;
  assign n1879 = ~g143 & n1149;
  assign n1880 = g143 & ~n1149;
  assign n1881 = ~n1158 & g157 & ~n1159;
  assign n1882 = ~g152 & n1876;
  assign n1161 = n1884 | n1897;
  assign n1884 = ~n806_1 & ~n1885;
  assign n1885 = ~n1886 & ~n1887;
  assign n1886 = ~g111 & n816_1;
  assign n1887 = g127 & ~n1888;
  assign n1888 = ~n1891 & ~g2584 & g119 & ~n1889;
  assign n1889 = ~n1161_1 & ~n1890 & ~n814 & ~n1143 & ~n813 & ~n815;
  assign n1890 = g89 & g107;
  assign n1891 = ~n1892 & ~n1896;
  assign n1892 = g697 & ~n1893;
  assign n1893 = ~n1894 & ~n1895;
  assign n1894 = g123 & ~n815;
  assign n1895 = ~n1143 & ~g123 & ~n1890 & ~n813;
  assign n1896 = ~g697 & n1893;
  assign n1897 = n806_1 & ~n1898;
  assign n1898 = ~n1901 & ~n823 & ~n1899 & ~n838;
  assign n1899 = ~n791_1 & ~n1192 & ~n1900;
  assign n1900 = n798 & n821_1 & ~g685 & ~g684;
  assign n1901 = ~n1902 & ~n963 & ~n1906;
  assign n1902 = ~n843 & ~n1903;
  assign n1903 = ~n1904 & ~n1905;
  assign n1904 = g293 & n791_1;
  assign n1905 = n797 & n861_1 & g688;
  assign n1906 = g658 & ~n1907;
  assign n1907 = ~n864 & n1746;
  assign n1166 = n1166_1 | n1909;
  assign n1909 = n1137 & ~n1910 & ~n1915;
  assign n1910 = g161 & ~n1911;
  assign n1911 = ~n1912 & ~n1913;
  assign n1912 = ~n1158 & g166 & ~n1159;
  assign n1913 = ~n1914 & ~n1158 & n1159 & ~n1878;
  assign n1914 = ~n1148 & ~n1154;
  assign n1915 = ~g161 & n1911;
  assign n1171 = n1917 | n1918;
  assign n1917 = g512 & ~n1329;
  assign n1918 = g693 & n1329;
  assign n1176 = n1920 | n1921;
  assign n1920 = g532 & ~n1022;
  assign n1921 = g690 & n1022;
  assign n1181 = n1055 | n1923;
  assign n1923 = n1028 & ~n1924 & ~n1931;
  assign n1924 = g64 & ~n1925;
  assign n1925 = ~n1926 & ~n1930;
  assign n1926 = ~n1047 & n1048 & ~n1927;
  assign n1927 = ~n1928 & ~n1929;
  assign n1928 = n1039 & ~g59 & ~g54 & n1038;
  assign n1929 = ~n1039 & g59 & g54 & n1043;
  assign n1930 = ~n1047 & g382 & ~n1048;
  assign n1931 = ~g64 & n1925;
  assign n1201 = n1055 | n1933;
  assign n1933 = n1028 & ~n1934 & ~n1941;
  assign n1934 = g59 & ~n1935;
  assign n1935 = ~n1936 & ~n1940;
  assign n1936 = ~n1047 & n1048 & ~n1937;
  assign n1937 = ~n1938 & ~n1939;
  assign n1938 = ~g54 & n1038 & n1039;
  assign n1939 = ~n1039 & g54 & n1043;
  assign n1940 = ~n1047 & g378 & ~n1048;
  assign n1941 = ~g59 & n1935;
  assign g3222 = g705;
  assign g3600 = g43;
  assign g4307 = g485;
  assign g4321 = g668;
  assign g4422 = g564;
  assign g5137 = g43;
  assign g5468 = g485;
  assign g5469 = g668;
  assign g5692 = 1'b0;
  assign g6282 = ~n713;
  assign g6728 = 1'b0;
  assign g1290 = g666;
  assign g4108 = g45;
  assign g4106 = g42;
  assign g4103 = g39;
  assign g1293 = g699;
  assign g4099 = g32;
  assign g4102 = g38;
  assign g4109 = g46;
  assign g4100 = g36;
  assign g4112 = g47;
  assign g4105 = g40;
  assign g4101 = g37;
  assign g4110 = g41;
  assign g4104 = g22;
  assign g4107 = g44;
  assign g4098 = g23;
  assign n151 = g2;
  assign n166 = ~n964;
  assign n171 = g18;
  assign n181 = g25;
  assign n186 = g571;
  assign n196 = g39;
  assign n201 = g29;
  assign n216 = g654;
  assign n221 = ~n1056_1;
  assign n236 = ~n1088;
  assign n266 = ~n742;
  assign n281 = g18;
  assign n316 = g646;
  assign n326 = g28;
  assign n336 = ~n1256;
  assign n341 = g650;
  assign n356 = g14;
  assign n366 = ~n1271;
  assign n381 = g634;
  assign n386 = g32;
  assign n401 = ~n1320;
  assign n406 = g28;
  assign n411 = ~n1216;
  assign n431 = g567;
  assign n456 = ~n1341;
  assign n481 = g10;
  assign n496 = ~g690;
  assign n501 = g664;
  assign n511 = g598;
  assign n531 = g567;
  assign n551 = ~g266;
  assign n576 = g663;
  assign n586 = ~n1423;
  assign n611 = g40;
  assign n626 = g1;
  assign n641 = g11;
  assign n646 = g37;
  assign n666 = g42;
  assign n691 = g24;
  assign n706 = g24;
  assign n721 = g654;
  assign n731 = g650;
  assign n736 = g7;
  assign n741 = g642;
  assign n761 = g6;
  assign n766 = g33;
  assign n771 = g38;
  assign n776 = ~n1415;
  assign n786 = g15;
  assign n791 = g19;
  assign n796 = g10;
  assign n811 = g45;
  assign n821 = ~n1360;
  assign n836 = g36;
  assign n841 = g606;
  assign n846 = g667;
  assign n861 = ~n1695;
  assign n866 = g42;
  assign n881 = ~n1708;
  assign n886 = g702;
  assign n891 = g665;
  assign n911 = g634;
  assign n916 = ~g691;
  assign n931 = g598;
  assign n936 = g646;
  assign n956 = ~n1746;
  assign n971 = ~n1474;
  assign n981 = g642;
  assign n991 = ~n1290;
  assign n1031 = g606;
  assign n1041 = ~n1790;
  assign n1051 = g46;
  assign n1066 = g571;
  assign n1091 = g1;
  assign n1101 = ~n910;
  assign n1106 = ~g47;
  assign n1151 = g6;
  assign n1156 = ~n1821;
  assign n1186 = g14;
  assign n1191 = g2;
  assign n1196 = g3;
  always @ (posedge clock) begin
    g678 <= n151;
    g332 <= n156;
    g123 <= n161;
    g207 <= n166;
    g695 <= n171;
    g461 <= n176;
    g18 <= n181;
    g292 <= n186;
    g331 <= n191;
    g689 <= n196;
    g24 <= n201;
    g465 <= n206;
    g84 <= n211;
    g291 <= n216;
    g676 <= n221;
    g622 <= n226;
    g117 <= n231;
    g278 <= n236;
    g128 <= n241;
    g598 <= n246;
    g554 <= n251;
    g496 <= n256;
    g179 <= n261;
    g48 <= n266;
    g590 <= n271;
    g551 <= n276;
    g682 <= n281;
    g11 <= n286;
    g606 <= n291;
    g188 <= n296;
    g646 <= n301;
    g327 <= n306;
    g361 <= n311;
    g289 <= n316;
    g398 <= n321;
    g684 <= n326;
    g619 <= n331;
    g208 <= n336;
    g248 <= n341;
    g390 <= n346;
    g625 <= n351;
    g681 <= n356;
    g437 <= n361;
    g276 <= n366;
    g3 <= n371;
    g323 <= n376;
    g224 <= n381;
    g685 <= n386;
    g43 <= n391;
    g157 <= n396;
    g282 <= n401;
    g697 <= n406;
    g206 <= n411;
    g449 <= n416;
    g118 <= n421;
    g528 <= n426;
    g284 <= n431;
    g426 <= n436;
    g634 <= n441;
    g669 <= n446;
    g520 <= n451;
    g281 <= n456;
    g175 <= n461;
    g15 <= n466;
    g631 <= n471;
    g69 <= n476;
    g693 <= n481;
    g337 <= n486;
    g457 <= n491;
    g486 <= n496;
    g471 <= n501;
    g328 <= n506;
    g285 <= n511;
    g418 <= n516;
    g402 <= n521;
    g297 <= n526;
    g212 <= n531;
    g410 <= n536;
    g430 <= n541;
    g33 <= n546;
    g662 <= n551;
    g453 <= n556;
    g269 <= n561;
    g574 <= n566;
    g441 <= n571;
    g664 <= n576;
    g349 <= n581;
    g211 <= n586;
    g586 <= n591;
    g571 <= n596;
    g29 <= n601;
    g326 <= n606;
    g698 <= n611;
    g654 <= n616;
    g293 <= n621;
    g690 <= n626;
    g445 <= n631;
    g374 <= n636;
    g6 <= n641;
    g687 <= n646;
    g357 <= n651;
    g386 <= n656;
    g504 <= n661;
    g665 <= n666;
    g166 <= n671;
    g541 <= n676;
    g74 <= n681;
    g338 <= n686;
    g696 <= n691;
    g516 <= n696;
    g536 <= n701;
    g683 <= n706;
    g353 <= n711;
    g545 <= n716;
    g254 <= n721;
    g341 <= n726;
    g290 <= n731;
    g2 <= n736;
    g287 <= n741;
    g336 <= n746;
    g345 <= n751;
    g628 <= n756;
    g679 <= n761;
    g28 <= n766;
    g688 <= n771;
    g283 <= n776;
    g613 <= n781;
    g10 <= n786;
    g14 <= n791;
    g680 <= n796;
    g143 <= n801;
    g672 <= n806;
    g667 <= n811;
    g366 <= n816;
    g279 <= n821;
    g492 <= n826;
    g170 <= n831;
    g686 <= n836;
    g288 <= n841;
    g638 <= n846;
    g602 <= n851;
    g642 <= n856;
    g280 <= n861;
    g663 <= n866;
    g610 <= n871;
    g148 <= n876;
    g209 <= n881;
    g675 <= n886;
    g478 <= n891;
    g122 <= n896;
    g54 <= n901;
    g594 <= n906;
    g286 <= n911;
    g489 <= n916;
    g616 <= n921;
    g79 <= n926;
    g218 <= n931;
    g242 <= n936;
    g578 <= n941;
    g184 <= n946;
    g119 <= n951;
    g668 <= n956;
    g139 <= n961;
    g422 <= n966;
    g210 <= n971;
    g394 <= n976;
    g230 <= n981;
    g25 <= n986;
    g204 <= n991;
    g658 <= n996;
    g650 <= n1001;
    g378 <= n1006;
    g508 <= n1011;
    g548 <= n1016;
    g370 <= n1021;
    g406 <= n1026;
    g236 <= n1031;
    g500 <= n1036;
    g205 <= n1041;
    g197 <= n1046;
    g666 <= n1051;
    g114 <= n1056;
    g524 <= n1061;
    g260 <= n1066;
    g111 <= n1071;
    g131 <= n1076;
    g7 <= n1081;
    g19 <= n1086;
    g677 <= n1091;
    g582 <= n1096;
    g485 <= n1101;
    g699 <= n1106;
    g193 <= n1111;
    g135 <= n1116;
    g382 <= n1121;
    g414 <= n1126;
    g434 <= n1131;
    g266 <= n1136;
    g49 <= n1141;
    g152 <= n1146;
    g692 <= n1151;
    g277 <= n1156;
    g127 <= n1161;
    g161 <= n1166;
    g512 <= n1171;
    g532 <= n1176;
    g64 <= n1181;
    g694 <= n1186;
    g691 <= n1191;
    g1 <= n1196;
    g59 <= n1201;
  end
endmodule


